module SimDualPortBRAM(
  input          clock,
  input          reset,
  input          io_web,
  input  [7:0]   io_addra,
  input  [7:0]   io_addrb,
  input  [127:0] io_dinb,
  output [127:0] io_douta
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [127:0] _RAND_14;
  reg [127:0] _RAND_15;
  reg [127:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [127:0] _RAND_19;
  reg [127:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [127:0] _RAND_22;
  reg [127:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [127:0] _RAND_25;
  reg [127:0] _RAND_26;
  reg [127:0] _RAND_27;
  reg [127:0] _RAND_28;
  reg [127:0] _RAND_29;
  reg [127:0] _RAND_30;
  reg [127:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [127:0] _RAND_33;
  reg [127:0] _RAND_34;
  reg [127:0] _RAND_35;
  reg [127:0] _RAND_36;
  reg [127:0] _RAND_37;
  reg [127:0] _RAND_38;
  reg [127:0] _RAND_39;
  reg [127:0] _RAND_40;
  reg [127:0] _RAND_41;
  reg [127:0] _RAND_42;
  reg [127:0] _RAND_43;
  reg [127:0] _RAND_44;
  reg [127:0] _RAND_45;
  reg [127:0] _RAND_46;
  reg [127:0] _RAND_47;
  reg [127:0] _RAND_48;
  reg [127:0] _RAND_49;
  reg [127:0] _RAND_50;
  reg [127:0] _RAND_51;
  reg [127:0] _RAND_52;
  reg [127:0] _RAND_53;
  reg [127:0] _RAND_54;
  reg [127:0] _RAND_55;
  reg [127:0] _RAND_56;
  reg [127:0] _RAND_57;
  reg [127:0] _RAND_58;
  reg [127:0] _RAND_59;
  reg [127:0] _RAND_60;
  reg [127:0] _RAND_61;
  reg [127:0] _RAND_62;
  reg [127:0] _RAND_63;
  reg [127:0] _RAND_64;
  reg [127:0] _RAND_65;
  reg [127:0] _RAND_66;
  reg [127:0] _RAND_67;
  reg [127:0] _RAND_68;
  reg [127:0] _RAND_69;
  reg [127:0] _RAND_70;
  reg [127:0] _RAND_71;
  reg [127:0] _RAND_72;
  reg [127:0] _RAND_73;
  reg [127:0] _RAND_74;
  reg [127:0] _RAND_75;
  reg [127:0] _RAND_76;
  reg [127:0] _RAND_77;
  reg [127:0] _RAND_78;
  reg [127:0] _RAND_79;
  reg [127:0] _RAND_80;
  reg [127:0] _RAND_81;
  reg [127:0] _RAND_82;
  reg [127:0] _RAND_83;
  reg [127:0] _RAND_84;
  reg [127:0] _RAND_85;
  reg [127:0] _RAND_86;
  reg [127:0] _RAND_87;
  reg [127:0] _RAND_88;
  reg [127:0] _RAND_89;
  reg [127:0] _RAND_90;
  reg [127:0] _RAND_91;
  reg [127:0] _RAND_92;
  reg [127:0] _RAND_93;
  reg [127:0] _RAND_94;
  reg [127:0] _RAND_95;
  reg [127:0] _RAND_96;
  reg [127:0] _RAND_97;
  reg [127:0] _RAND_98;
  reg [127:0] _RAND_99;
  reg [127:0] _RAND_100;
  reg [127:0] _RAND_101;
  reg [127:0] _RAND_102;
  reg [127:0] _RAND_103;
  reg [127:0] _RAND_104;
  reg [127:0] _RAND_105;
  reg [127:0] _RAND_106;
  reg [127:0] _RAND_107;
  reg [127:0] _RAND_108;
  reg [127:0] _RAND_109;
  reg [127:0] _RAND_110;
  reg [127:0] _RAND_111;
  reg [127:0] _RAND_112;
  reg [127:0] _RAND_113;
  reg [127:0] _RAND_114;
  reg [127:0] _RAND_115;
  reg [127:0] _RAND_116;
  reg [127:0] _RAND_117;
  reg [127:0] _RAND_118;
  reg [127:0] _RAND_119;
  reg [127:0] _RAND_120;
  reg [127:0] _RAND_121;
  reg [127:0] _RAND_122;
  reg [127:0] _RAND_123;
  reg [127:0] _RAND_124;
  reg [127:0] _RAND_125;
  reg [127:0] _RAND_126;
  reg [127:0] _RAND_127;
  reg [127:0] _RAND_128;
  reg [127:0] _RAND_129;
  reg [127:0] _RAND_130;
  reg [127:0] _RAND_131;
  reg [127:0] _RAND_132;
  reg [127:0] _RAND_133;
  reg [127:0] _RAND_134;
  reg [127:0] _RAND_135;
  reg [127:0] _RAND_136;
  reg [127:0] _RAND_137;
  reg [127:0] _RAND_138;
  reg [127:0] _RAND_139;
  reg [127:0] _RAND_140;
  reg [127:0] _RAND_141;
  reg [127:0] _RAND_142;
  reg [127:0] _RAND_143;
  reg [127:0] _RAND_144;
  reg [127:0] _RAND_145;
  reg [127:0] _RAND_146;
  reg [127:0] _RAND_147;
  reg [127:0] _RAND_148;
  reg [127:0] _RAND_149;
  reg [127:0] _RAND_150;
  reg [127:0] _RAND_151;
  reg [127:0] _RAND_152;
  reg [127:0] _RAND_153;
  reg [127:0] _RAND_154;
  reg [127:0] _RAND_155;
  reg [127:0] _RAND_156;
  reg [127:0] _RAND_157;
  reg [127:0] _RAND_158;
  reg [127:0] _RAND_159;
  reg [127:0] _RAND_160;
  reg [127:0] _RAND_161;
  reg [127:0] _RAND_162;
  reg [127:0] _RAND_163;
  reg [127:0] _RAND_164;
  reg [127:0] _RAND_165;
  reg [127:0] _RAND_166;
  reg [127:0] _RAND_167;
  reg [127:0] _RAND_168;
  reg [127:0] _RAND_169;
  reg [127:0] _RAND_170;
  reg [127:0] _RAND_171;
  reg [127:0] _RAND_172;
  reg [127:0] _RAND_173;
  reg [127:0] _RAND_174;
  reg [127:0] _RAND_175;
  reg [127:0] _RAND_176;
  reg [127:0] _RAND_177;
  reg [127:0] _RAND_178;
  reg [127:0] _RAND_179;
  reg [127:0] _RAND_180;
  reg [127:0] _RAND_181;
  reg [127:0] _RAND_182;
  reg [127:0] _RAND_183;
  reg [127:0] _RAND_184;
  reg [127:0] _RAND_185;
  reg [127:0] _RAND_186;
  reg [127:0] _RAND_187;
  reg [127:0] _RAND_188;
  reg [127:0] _RAND_189;
  reg [127:0] _RAND_190;
  reg [127:0] _RAND_191;
  reg [127:0] _RAND_192;
  reg [127:0] _RAND_193;
  reg [127:0] _RAND_194;
  reg [127:0] _RAND_195;
  reg [127:0] _RAND_196;
  reg [127:0] _RAND_197;
  reg [127:0] _RAND_198;
  reg [127:0] _RAND_199;
  reg [127:0] _RAND_200;
  reg [127:0] _RAND_201;
  reg [127:0] _RAND_202;
  reg [127:0] _RAND_203;
  reg [127:0] _RAND_204;
  reg [127:0] _RAND_205;
  reg [127:0] _RAND_206;
  reg [127:0] _RAND_207;
  reg [127:0] _RAND_208;
  reg [127:0] _RAND_209;
  reg [127:0] _RAND_210;
  reg [127:0] _RAND_211;
  reg [127:0] _RAND_212;
  reg [127:0] _RAND_213;
  reg [127:0] _RAND_214;
  reg [127:0] _RAND_215;
  reg [127:0] _RAND_216;
  reg [127:0] _RAND_217;
  reg [127:0] _RAND_218;
  reg [127:0] _RAND_219;
  reg [127:0] _RAND_220;
  reg [127:0] _RAND_221;
  reg [127:0] _RAND_222;
  reg [127:0] _RAND_223;
  reg [127:0] _RAND_224;
  reg [127:0] _RAND_225;
  reg [127:0] _RAND_226;
  reg [127:0] _RAND_227;
  reg [127:0] _RAND_228;
  reg [127:0] _RAND_229;
  reg [127:0] _RAND_230;
  reg [127:0] _RAND_231;
  reg [127:0] _RAND_232;
  reg [127:0] _RAND_233;
  reg [127:0] _RAND_234;
  reg [127:0] _RAND_235;
  reg [127:0] _RAND_236;
  reg [127:0] _RAND_237;
  reg [127:0] _RAND_238;
  reg [127:0] _RAND_239;
  reg [127:0] _RAND_240;
  reg [127:0] _RAND_241;
  reg [127:0] _RAND_242;
  reg [127:0] _RAND_243;
  reg [127:0] _RAND_244;
  reg [127:0] _RAND_245;
  reg [127:0] _RAND_246;
  reg [127:0] _RAND_247;
  reg [127:0] _RAND_248;
  reg [127:0] _RAND_249;
  reg [127:0] _RAND_250;
  reg [127:0] _RAND_251;
  reg [127:0] _RAND_252;
  reg [127:0] _RAND_253;
  reg [127:0] _RAND_254;
  reg [127:0] _RAND_255;
  reg [127:0] _RAND_256;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] mem_0; // @[RAM.scala 41:22]
  reg [127:0] mem_1; // @[RAM.scala 41:22]
  reg [127:0] mem_2; // @[RAM.scala 41:22]
  reg [127:0] mem_3; // @[RAM.scala 41:22]
  reg [127:0] mem_4; // @[RAM.scala 41:22]
  reg [127:0] mem_5; // @[RAM.scala 41:22]
  reg [127:0] mem_6; // @[RAM.scala 41:22]
  reg [127:0] mem_7; // @[RAM.scala 41:22]
  reg [127:0] mem_8; // @[RAM.scala 41:22]
  reg [127:0] mem_9; // @[RAM.scala 41:22]
  reg [127:0] mem_10; // @[RAM.scala 41:22]
  reg [127:0] mem_11; // @[RAM.scala 41:22]
  reg [127:0] mem_12; // @[RAM.scala 41:22]
  reg [127:0] mem_13; // @[RAM.scala 41:22]
  reg [127:0] mem_14; // @[RAM.scala 41:22]
  reg [127:0] mem_15; // @[RAM.scala 41:22]
  reg [127:0] mem_16; // @[RAM.scala 41:22]
  reg [127:0] mem_17; // @[RAM.scala 41:22]
  reg [127:0] mem_18; // @[RAM.scala 41:22]
  reg [127:0] mem_19; // @[RAM.scala 41:22]
  reg [127:0] mem_20; // @[RAM.scala 41:22]
  reg [127:0] mem_21; // @[RAM.scala 41:22]
  reg [127:0] mem_22; // @[RAM.scala 41:22]
  reg [127:0] mem_23; // @[RAM.scala 41:22]
  reg [127:0] mem_24; // @[RAM.scala 41:22]
  reg [127:0] mem_25; // @[RAM.scala 41:22]
  reg [127:0] mem_26; // @[RAM.scala 41:22]
  reg [127:0] mem_27; // @[RAM.scala 41:22]
  reg [127:0] mem_28; // @[RAM.scala 41:22]
  reg [127:0] mem_29; // @[RAM.scala 41:22]
  reg [127:0] mem_30; // @[RAM.scala 41:22]
  reg [127:0] mem_31; // @[RAM.scala 41:22]
  reg [127:0] mem_32; // @[RAM.scala 41:22]
  reg [127:0] mem_33; // @[RAM.scala 41:22]
  reg [127:0] mem_34; // @[RAM.scala 41:22]
  reg [127:0] mem_35; // @[RAM.scala 41:22]
  reg [127:0] mem_36; // @[RAM.scala 41:22]
  reg [127:0] mem_37; // @[RAM.scala 41:22]
  reg [127:0] mem_38; // @[RAM.scala 41:22]
  reg [127:0] mem_39; // @[RAM.scala 41:22]
  reg [127:0] mem_40; // @[RAM.scala 41:22]
  reg [127:0] mem_41; // @[RAM.scala 41:22]
  reg [127:0] mem_42; // @[RAM.scala 41:22]
  reg [127:0] mem_43; // @[RAM.scala 41:22]
  reg [127:0] mem_44; // @[RAM.scala 41:22]
  reg [127:0] mem_45; // @[RAM.scala 41:22]
  reg [127:0] mem_46; // @[RAM.scala 41:22]
  reg [127:0] mem_47; // @[RAM.scala 41:22]
  reg [127:0] mem_48; // @[RAM.scala 41:22]
  reg [127:0] mem_49; // @[RAM.scala 41:22]
  reg [127:0] mem_50; // @[RAM.scala 41:22]
  reg [127:0] mem_51; // @[RAM.scala 41:22]
  reg [127:0] mem_52; // @[RAM.scala 41:22]
  reg [127:0] mem_53; // @[RAM.scala 41:22]
  reg [127:0] mem_54; // @[RAM.scala 41:22]
  reg [127:0] mem_55; // @[RAM.scala 41:22]
  reg [127:0] mem_56; // @[RAM.scala 41:22]
  reg [127:0] mem_57; // @[RAM.scala 41:22]
  reg [127:0] mem_58; // @[RAM.scala 41:22]
  reg [127:0] mem_59; // @[RAM.scala 41:22]
  reg [127:0] mem_60; // @[RAM.scala 41:22]
  reg [127:0] mem_61; // @[RAM.scala 41:22]
  reg [127:0] mem_62; // @[RAM.scala 41:22]
  reg [127:0] mem_63; // @[RAM.scala 41:22]
  reg [127:0] mem_64; // @[RAM.scala 41:22]
  reg [127:0] mem_65; // @[RAM.scala 41:22]
  reg [127:0] mem_66; // @[RAM.scala 41:22]
  reg [127:0] mem_67; // @[RAM.scala 41:22]
  reg [127:0] mem_68; // @[RAM.scala 41:22]
  reg [127:0] mem_69; // @[RAM.scala 41:22]
  reg [127:0] mem_70; // @[RAM.scala 41:22]
  reg [127:0] mem_71; // @[RAM.scala 41:22]
  reg [127:0] mem_72; // @[RAM.scala 41:22]
  reg [127:0] mem_73; // @[RAM.scala 41:22]
  reg [127:0] mem_74; // @[RAM.scala 41:22]
  reg [127:0] mem_75; // @[RAM.scala 41:22]
  reg [127:0] mem_76; // @[RAM.scala 41:22]
  reg [127:0] mem_77; // @[RAM.scala 41:22]
  reg [127:0] mem_78; // @[RAM.scala 41:22]
  reg [127:0] mem_79; // @[RAM.scala 41:22]
  reg [127:0] mem_80; // @[RAM.scala 41:22]
  reg [127:0] mem_81; // @[RAM.scala 41:22]
  reg [127:0] mem_82; // @[RAM.scala 41:22]
  reg [127:0] mem_83; // @[RAM.scala 41:22]
  reg [127:0] mem_84; // @[RAM.scala 41:22]
  reg [127:0] mem_85; // @[RAM.scala 41:22]
  reg [127:0] mem_86; // @[RAM.scala 41:22]
  reg [127:0] mem_87; // @[RAM.scala 41:22]
  reg [127:0] mem_88; // @[RAM.scala 41:22]
  reg [127:0] mem_89; // @[RAM.scala 41:22]
  reg [127:0] mem_90; // @[RAM.scala 41:22]
  reg [127:0] mem_91; // @[RAM.scala 41:22]
  reg [127:0] mem_92; // @[RAM.scala 41:22]
  reg [127:0] mem_93; // @[RAM.scala 41:22]
  reg [127:0] mem_94; // @[RAM.scala 41:22]
  reg [127:0] mem_95; // @[RAM.scala 41:22]
  reg [127:0] mem_96; // @[RAM.scala 41:22]
  reg [127:0] mem_97; // @[RAM.scala 41:22]
  reg [127:0] mem_98; // @[RAM.scala 41:22]
  reg [127:0] mem_99; // @[RAM.scala 41:22]
  reg [127:0] mem_100; // @[RAM.scala 41:22]
  reg [127:0] mem_101; // @[RAM.scala 41:22]
  reg [127:0] mem_102; // @[RAM.scala 41:22]
  reg [127:0] mem_103; // @[RAM.scala 41:22]
  reg [127:0] mem_104; // @[RAM.scala 41:22]
  reg [127:0] mem_105; // @[RAM.scala 41:22]
  reg [127:0] mem_106; // @[RAM.scala 41:22]
  reg [127:0] mem_107; // @[RAM.scala 41:22]
  reg [127:0] mem_108; // @[RAM.scala 41:22]
  reg [127:0] mem_109; // @[RAM.scala 41:22]
  reg [127:0] mem_110; // @[RAM.scala 41:22]
  reg [127:0] mem_111; // @[RAM.scala 41:22]
  reg [127:0] mem_112; // @[RAM.scala 41:22]
  reg [127:0] mem_113; // @[RAM.scala 41:22]
  reg [127:0] mem_114; // @[RAM.scala 41:22]
  reg [127:0] mem_115; // @[RAM.scala 41:22]
  reg [127:0] mem_116; // @[RAM.scala 41:22]
  reg [127:0] mem_117; // @[RAM.scala 41:22]
  reg [127:0] mem_118; // @[RAM.scala 41:22]
  reg [127:0] mem_119; // @[RAM.scala 41:22]
  reg [127:0] mem_120; // @[RAM.scala 41:22]
  reg [127:0] mem_121; // @[RAM.scala 41:22]
  reg [127:0] mem_122; // @[RAM.scala 41:22]
  reg [127:0] mem_123; // @[RAM.scala 41:22]
  reg [127:0] mem_124; // @[RAM.scala 41:22]
  reg [127:0] mem_125; // @[RAM.scala 41:22]
  reg [127:0] mem_126; // @[RAM.scala 41:22]
  reg [127:0] mem_127; // @[RAM.scala 41:22]
  reg [127:0] mem_128; // @[RAM.scala 41:22]
  reg [127:0] mem_129; // @[RAM.scala 41:22]
  reg [127:0] mem_130; // @[RAM.scala 41:22]
  reg [127:0] mem_131; // @[RAM.scala 41:22]
  reg [127:0] mem_132; // @[RAM.scala 41:22]
  reg [127:0] mem_133; // @[RAM.scala 41:22]
  reg [127:0] mem_134; // @[RAM.scala 41:22]
  reg [127:0] mem_135; // @[RAM.scala 41:22]
  reg [127:0] mem_136; // @[RAM.scala 41:22]
  reg [127:0] mem_137; // @[RAM.scala 41:22]
  reg [127:0] mem_138; // @[RAM.scala 41:22]
  reg [127:0] mem_139; // @[RAM.scala 41:22]
  reg [127:0] mem_140; // @[RAM.scala 41:22]
  reg [127:0] mem_141; // @[RAM.scala 41:22]
  reg [127:0] mem_142; // @[RAM.scala 41:22]
  reg [127:0] mem_143; // @[RAM.scala 41:22]
  reg [127:0] mem_144; // @[RAM.scala 41:22]
  reg [127:0] mem_145; // @[RAM.scala 41:22]
  reg [127:0] mem_146; // @[RAM.scala 41:22]
  reg [127:0] mem_147; // @[RAM.scala 41:22]
  reg [127:0] mem_148; // @[RAM.scala 41:22]
  reg [127:0] mem_149; // @[RAM.scala 41:22]
  reg [127:0] mem_150; // @[RAM.scala 41:22]
  reg [127:0] mem_151; // @[RAM.scala 41:22]
  reg [127:0] mem_152; // @[RAM.scala 41:22]
  reg [127:0] mem_153; // @[RAM.scala 41:22]
  reg [127:0] mem_154; // @[RAM.scala 41:22]
  reg [127:0] mem_155; // @[RAM.scala 41:22]
  reg [127:0] mem_156; // @[RAM.scala 41:22]
  reg [127:0] mem_157; // @[RAM.scala 41:22]
  reg [127:0] mem_158; // @[RAM.scala 41:22]
  reg [127:0] mem_159; // @[RAM.scala 41:22]
  reg [127:0] mem_160; // @[RAM.scala 41:22]
  reg [127:0] mem_161; // @[RAM.scala 41:22]
  reg [127:0] mem_162; // @[RAM.scala 41:22]
  reg [127:0] mem_163; // @[RAM.scala 41:22]
  reg [127:0] mem_164; // @[RAM.scala 41:22]
  reg [127:0] mem_165; // @[RAM.scala 41:22]
  reg [127:0] mem_166; // @[RAM.scala 41:22]
  reg [127:0] mem_167; // @[RAM.scala 41:22]
  reg [127:0] mem_168; // @[RAM.scala 41:22]
  reg [127:0] mem_169; // @[RAM.scala 41:22]
  reg [127:0] mem_170; // @[RAM.scala 41:22]
  reg [127:0] mem_171; // @[RAM.scala 41:22]
  reg [127:0] mem_172; // @[RAM.scala 41:22]
  reg [127:0] mem_173; // @[RAM.scala 41:22]
  reg [127:0] mem_174; // @[RAM.scala 41:22]
  reg [127:0] mem_175; // @[RAM.scala 41:22]
  reg [127:0] mem_176; // @[RAM.scala 41:22]
  reg [127:0] mem_177; // @[RAM.scala 41:22]
  reg [127:0] mem_178; // @[RAM.scala 41:22]
  reg [127:0] mem_179; // @[RAM.scala 41:22]
  reg [127:0] mem_180; // @[RAM.scala 41:22]
  reg [127:0] mem_181; // @[RAM.scala 41:22]
  reg [127:0] mem_182; // @[RAM.scala 41:22]
  reg [127:0] mem_183; // @[RAM.scala 41:22]
  reg [127:0] mem_184; // @[RAM.scala 41:22]
  reg [127:0] mem_185; // @[RAM.scala 41:22]
  reg [127:0] mem_186; // @[RAM.scala 41:22]
  reg [127:0] mem_187; // @[RAM.scala 41:22]
  reg [127:0] mem_188; // @[RAM.scala 41:22]
  reg [127:0] mem_189; // @[RAM.scala 41:22]
  reg [127:0] mem_190; // @[RAM.scala 41:22]
  reg [127:0] mem_191; // @[RAM.scala 41:22]
  reg [127:0] mem_192; // @[RAM.scala 41:22]
  reg [127:0] mem_193; // @[RAM.scala 41:22]
  reg [127:0] mem_194; // @[RAM.scala 41:22]
  reg [127:0] mem_195; // @[RAM.scala 41:22]
  reg [127:0] mem_196; // @[RAM.scala 41:22]
  reg [127:0] mem_197; // @[RAM.scala 41:22]
  reg [127:0] mem_198; // @[RAM.scala 41:22]
  reg [127:0] mem_199; // @[RAM.scala 41:22]
  reg [127:0] mem_200; // @[RAM.scala 41:22]
  reg [127:0] mem_201; // @[RAM.scala 41:22]
  reg [127:0] mem_202; // @[RAM.scala 41:22]
  reg [127:0] mem_203; // @[RAM.scala 41:22]
  reg [127:0] mem_204; // @[RAM.scala 41:22]
  reg [127:0] mem_205; // @[RAM.scala 41:22]
  reg [127:0] mem_206; // @[RAM.scala 41:22]
  reg [127:0] mem_207; // @[RAM.scala 41:22]
  reg [127:0] mem_208; // @[RAM.scala 41:22]
  reg [127:0] mem_209; // @[RAM.scala 41:22]
  reg [127:0] mem_210; // @[RAM.scala 41:22]
  reg [127:0] mem_211; // @[RAM.scala 41:22]
  reg [127:0] mem_212; // @[RAM.scala 41:22]
  reg [127:0] mem_213; // @[RAM.scala 41:22]
  reg [127:0] mem_214; // @[RAM.scala 41:22]
  reg [127:0] mem_215; // @[RAM.scala 41:22]
  reg [127:0] mem_216; // @[RAM.scala 41:22]
  reg [127:0] mem_217; // @[RAM.scala 41:22]
  reg [127:0] mem_218; // @[RAM.scala 41:22]
  reg [127:0] mem_219; // @[RAM.scala 41:22]
  reg [127:0] mem_220; // @[RAM.scala 41:22]
  reg [127:0] mem_221; // @[RAM.scala 41:22]
  reg [127:0] mem_222; // @[RAM.scala 41:22]
  reg [127:0] mem_223; // @[RAM.scala 41:22]
  reg [127:0] mem_224; // @[RAM.scala 41:22]
  reg [127:0] mem_225; // @[RAM.scala 41:22]
  reg [127:0] mem_226; // @[RAM.scala 41:22]
  reg [127:0] mem_227; // @[RAM.scala 41:22]
  reg [127:0] mem_228; // @[RAM.scala 41:22]
  reg [127:0] mem_229; // @[RAM.scala 41:22]
  reg [127:0] mem_230; // @[RAM.scala 41:22]
  reg [127:0] mem_231; // @[RAM.scala 41:22]
  reg [127:0] mem_232; // @[RAM.scala 41:22]
  reg [127:0] mem_233; // @[RAM.scala 41:22]
  reg [127:0] mem_234; // @[RAM.scala 41:22]
  reg [127:0] mem_235; // @[RAM.scala 41:22]
  reg [127:0] mem_236; // @[RAM.scala 41:22]
  reg [127:0] mem_237; // @[RAM.scala 41:22]
  reg [127:0] mem_238; // @[RAM.scala 41:22]
  reg [127:0] mem_239; // @[RAM.scala 41:22]
  reg [127:0] mem_240; // @[RAM.scala 41:22]
  reg [127:0] mem_241; // @[RAM.scala 41:22]
  reg [127:0] mem_242; // @[RAM.scala 41:22]
  reg [127:0] mem_243; // @[RAM.scala 41:22]
  reg [127:0] mem_244; // @[RAM.scala 41:22]
  reg [127:0] mem_245; // @[RAM.scala 41:22]
  reg [127:0] mem_246; // @[RAM.scala 41:22]
  reg [127:0] mem_247; // @[RAM.scala 41:22]
  reg [127:0] mem_248; // @[RAM.scala 41:22]
  reg [127:0] mem_249; // @[RAM.scala 41:22]
  reg [127:0] mem_250; // @[RAM.scala 41:22]
  reg [127:0] mem_251; // @[RAM.scala 41:22]
  reg [127:0] mem_252; // @[RAM.scala 41:22]
  reg [127:0] mem_253; // @[RAM.scala 41:22]
  reg [127:0] mem_254; // @[RAM.scala 41:22]
  reg [127:0] mem_255; // @[RAM.scala 41:22]
  reg [127:0] io_douta_REG; // @[RAM.scala 43:24]
  wire [127:0] _GEN_1 = 8'h1 == io_addra ? mem_1 : mem_0; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_2 = 8'h2 == io_addra ? mem_2 : _GEN_1; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_3 = 8'h3 == io_addra ? mem_3 : _GEN_2; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_4 = 8'h4 == io_addra ? mem_4 : _GEN_3; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_5 = 8'h5 == io_addra ? mem_5 : _GEN_4; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_6 = 8'h6 == io_addra ? mem_6 : _GEN_5; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_7 = 8'h7 == io_addra ? mem_7 : _GEN_6; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_8 = 8'h8 == io_addra ? mem_8 : _GEN_7; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_9 = 8'h9 == io_addra ? mem_9 : _GEN_8; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_10 = 8'ha == io_addra ? mem_10 : _GEN_9; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_11 = 8'hb == io_addra ? mem_11 : _GEN_10; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_12 = 8'hc == io_addra ? mem_12 : _GEN_11; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_13 = 8'hd == io_addra ? mem_13 : _GEN_12; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_14 = 8'he == io_addra ? mem_14 : _GEN_13; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_15 = 8'hf == io_addra ? mem_15 : _GEN_14; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_16 = 8'h10 == io_addra ? mem_16 : _GEN_15; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_17 = 8'h11 == io_addra ? mem_17 : _GEN_16; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_18 = 8'h12 == io_addra ? mem_18 : _GEN_17; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_19 = 8'h13 == io_addra ? mem_19 : _GEN_18; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_20 = 8'h14 == io_addra ? mem_20 : _GEN_19; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_21 = 8'h15 == io_addra ? mem_21 : _GEN_20; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_22 = 8'h16 == io_addra ? mem_22 : _GEN_21; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_23 = 8'h17 == io_addra ? mem_23 : _GEN_22; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_24 = 8'h18 == io_addra ? mem_24 : _GEN_23; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_25 = 8'h19 == io_addra ? mem_25 : _GEN_24; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_26 = 8'h1a == io_addra ? mem_26 : _GEN_25; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_27 = 8'h1b == io_addra ? mem_27 : _GEN_26; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_28 = 8'h1c == io_addra ? mem_28 : _GEN_27; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_29 = 8'h1d == io_addra ? mem_29 : _GEN_28; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_30 = 8'h1e == io_addra ? mem_30 : _GEN_29; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_31 = 8'h1f == io_addra ? mem_31 : _GEN_30; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_32 = 8'h20 == io_addra ? mem_32 : _GEN_31; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_33 = 8'h21 == io_addra ? mem_33 : _GEN_32; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_34 = 8'h22 == io_addra ? mem_34 : _GEN_33; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_35 = 8'h23 == io_addra ? mem_35 : _GEN_34; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_36 = 8'h24 == io_addra ? mem_36 : _GEN_35; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_37 = 8'h25 == io_addra ? mem_37 : _GEN_36; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_38 = 8'h26 == io_addra ? mem_38 : _GEN_37; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_39 = 8'h27 == io_addra ? mem_39 : _GEN_38; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_40 = 8'h28 == io_addra ? mem_40 : _GEN_39; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_41 = 8'h29 == io_addra ? mem_41 : _GEN_40; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_42 = 8'h2a == io_addra ? mem_42 : _GEN_41; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_43 = 8'h2b == io_addra ? mem_43 : _GEN_42; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_44 = 8'h2c == io_addra ? mem_44 : _GEN_43; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_45 = 8'h2d == io_addra ? mem_45 : _GEN_44; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_46 = 8'h2e == io_addra ? mem_46 : _GEN_45; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_47 = 8'h2f == io_addra ? mem_47 : _GEN_46; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_48 = 8'h30 == io_addra ? mem_48 : _GEN_47; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_49 = 8'h31 == io_addra ? mem_49 : _GEN_48; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_50 = 8'h32 == io_addra ? mem_50 : _GEN_49; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_51 = 8'h33 == io_addra ? mem_51 : _GEN_50; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_52 = 8'h34 == io_addra ? mem_52 : _GEN_51; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_53 = 8'h35 == io_addra ? mem_53 : _GEN_52; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_54 = 8'h36 == io_addra ? mem_54 : _GEN_53; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_55 = 8'h37 == io_addra ? mem_55 : _GEN_54; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_56 = 8'h38 == io_addra ? mem_56 : _GEN_55; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_57 = 8'h39 == io_addra ? mem_57 : _GEN_56; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_58 = 8'h3a == io_addra ? mem_58 : _GEN_57; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_59 = 8'h3b == io_addra ? mem_59 : _GEN_58; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_60 = 8'h3c == io_addra ? mem_60 : _GEN_59; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_61 = 8'h3d == io_addra ? mem_61 : _GEN_60; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_62 = 8'h3e == io_addra ? mem_62 : _GEN_61; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_63 = 8'h3f == io_addra ? mem_63 : _GEN_62; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_64 = 8'h40 == io_addra ? mem_64 : _GEN_63; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_65 = 8'h41 == io_addra ? mem_65 : _GEN_64; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_66 = 8'h42 == io_addra ? mem_66 : _GEN_65; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_67 = 8'h43 == io_addra ? mem_67 : _GEN_66; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_68 = 8'h44 == io_addra ? mem_68 : _GEN_67; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_69 = 8'h45 == io_addra ? mem_69 : _GEN_68; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_70 = 8'h46 == io_addra ? mem_70 : _GEN_69; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_71 = 8'h47 == io_addra ? mem_71 : _GEN_70; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_72 = 8'h48 == io_addra ? mem_72 : _GEN_71; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_73 = 8'h49 == io_addra ? mem_73 : _GEN_72; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_74 = 8'h4a == io_addra ? mem_74 : _GEN_73; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_75 = 8'h4b == io_addra ? mem_75 : _GEN_74; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_76 = 8'h4c == io_addra ? mem_76 : _GEN_75; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_77 = 8'h4d == io_addra ? mem_77 : _GEN_76; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_78 = 8'h4e == io_addra ? mem_78 : _GEN_77; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_79 = 8'h4f == io_addra ? mem_79 : _GEN_78; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_80 = 8'h50 == io_addra ? mem_80 : _GEN_79; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_81 = 8'h51 == io_addra ? mem_81 : _GEN_80; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_82 = 8'h52 == io_addra ? mem_82 : _GEN_81; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_83 = 8'h53 == io_addra ? mem_83 : _GEN_82; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_84 = 8'h54 == io_addra ? mem_84 : _GEN_83; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_85 = 8'h55 == io_addra ? mem_85 : _GEN_84; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_86 = 8'h56 == io_addra ? mem_86 : _GEN_85; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_87 = 8'h57 == io_addra ? mem_87 : _GEN_86; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_88 = 8'h58 == io_addra ? mem_88 : _GEN_87; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_89 = 8'h59 == io_addra ? mem_89 : _GEN_88; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_90 = 8'h5a == io_addra ? mem_90 : _GEN_89; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_91 = 8'h5b == io_addra ? mem_91 : _GEN_90; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_92 = 8'h5c == io_addra ? mem_92 : _GEN_91; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_93 = 8'h5d == io_addra ? mem_93 : _GEN_92; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_94 = 8'h5e == io_addra ? mem_94 : _GEN_93; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_95 = 8'h5f == io_addra ? mem_95 : _GEN_94; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_96 = 8'h60 == io_addra ? mem_96 : _GEN_95; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_97 = 8'h61 == io_addra ? mem_97 : _GEN_96; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_98 = 8'h62 == io_addra ? mem_98 : _GEN_97; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_99 = 8'h63 == io_addra ? mem_99 : _GEN_98; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_100 = 8'h64 == io_addra ? mem_100 : _GEN_99; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_101 = 8'h65 == io_addra ? mem_101 : _GEN_100; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_102 = 8'h66 == io_addra ? mem_102 : _GEN_101; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_103 = 8'h67 == io_addra ? mem_103 : _GEN_102; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_104 = 8'h68 == io_addra ? mem_104 : _GEN_103; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_105 = 8'h69 == io_addra ? mem_105 : _GEN_104; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_106 = 8'h6a == io_addra ? mem_106 : _GEN_105; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_107 = 8'h6b == io_addra ? mem_107 : _GEN_106; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_108 = 8'h6c == io_addra ? mem_108 : _GEN_107; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_109 = 8'h6d == io_addra ? mem_109 : _GEN_108; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_110 = 8'h6e == io_addra ? mem_110 : _GEN_109; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_111 = 8'h6f == io_addra ? mem_111 : _GEN_110; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_112 = 8'h70 == io_addra ? mem_112 : _GEN_111; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_113 = 8'h71 == io_addra ? mem_113 : _GEN_112; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_114 = 8'h72 == io_addra ? mem_114 : _GEN_113; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_115 = 8'h73 == io_addra ? mem_115 : _GEN_114; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_116 = 8'h74 == io_addra ? mem_116 : _GEN_115; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_117 = 8'h75 == io_addra ? mem_117 : _GEN_116; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_118 = 8'h76 == io_addra ? mem_118 : _GEN_117; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_119 = 8'h77 == io_addra ? mem_119 : _GEN_118; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_120 = 8'h78 == io_addra ? mem_120 : _GEN_119; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_121 = 8'h79 == io_addra ? mem_121 : _GEN_120; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_122 = 8'h7a == io_addra ? mem_122 : _GEN_121; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_123 = 8'h7b == io_addra ? mem_123 : _GEN_122; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_124 = 8'h7c == io_addra ? mem_124 : _GEN_123; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_125 = 8'h7d == io_addra ? mem_125 : _GEN_124; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_126 = 8'h7e == io_addra ? mem_126 : _GEN_125; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_127 = 8'h7f == io_addra ? mem_127 : _GEN_126; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_128 = 8'h80 == io_addra ? mem_128 : _GEN_127; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_129 = 8'h81 == io_addra ? mem_129 : _GEN_128; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_130 = 8'h82 == io_addra ? mem_130 : _GEN_129; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_131 = 8'h83 == io_addra ? mem_131 : _GEN_130; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_132 = 8'h84 == io_addra ? mem_132 : _GEN_131; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_133 = 8'h85 == io_addra ? mem_133 : _GEN_132; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_134 = 8'h86 == io_addra ? mem_134 : _GEN_133; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_135 = 8'h87 == io_addra ? mem_135 : _GEN_134; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_136 = 8'h88 == io_addra ? mem_136 : _GEN_135; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_137 = 8'h89 == io_addra ? mem_137 : _GEN_136; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_138 = 8'h8a == io_addra ? mem_138 : _GEN_137; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_139 = 8'h8b == io_addra ? mem_139 : _GEN_138; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_140 = 8'h8c == io_addra ? mem_140 : _GEN_139; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_141 = 8'h8d == io_addra ? mem_141 : _GEN_140; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_142 = 8'h8e == io_addra ? mem_142 : _GEN_141; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_143 = 8'h8f == io_addra ? mem_143 : _GEN_142; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_144 = 8'h90 == io_addra ? mem_144 : _GEN_143; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_145 = 8'h91 == io_addra ? mem_145 : _GEN_144; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_146 = 8'h92 == io_addra ? mem_146 : _GEN_145; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_147 = 8'h93 == io_addra ? mem_147 : _GEN_146; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_148 = 8'h94 == io_addra ? mem_148 : _GEN_147; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_149 = 8'h95 == io_addra ? mem_149 : _GEN_148; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_150 = 8'h96 == io_addra ? mem_150 : _GEN_149; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_151 = 8'h97 == io_addra ? mem_151 : _GEN_150; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_152 = 8'h98 == io_addra ? mem_152 : _GEN_151; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_153 = 8'h99 == io_addra ? mem_153 : _GEN_152; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_154 = 8'h9a == io_addra ? mem_154 : _GEN_153; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_155 = 8'h9b == io_addra ? mem_155 : _GEN_154; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_156 = 8'h9c == io_addra ? mem_156 : _GEN_155; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_157 = 8'h9d == io_addra ? mem_157 : _GEN_156; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_158 = 8'h9e == io_addra ? mem_158 : _GEN_157; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_159 = 8'h9f == io_addra ? mem_159 : _GEN_158; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_160 = 8'ha0 == io_addra ? mem_160 : _GEN_159; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_161 = 8'ha1 == io_addra ? mem_161 : _GEN_160; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_162 = 8'ha2 == io_addra ? mem_162 : _GEN_161; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_163 = 8'ha3 == io_addra ? mem_163 : _GEN_162; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_164 = 8'ha4 == io_addra ? mem_164 : _GEN_163; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_165 = 8'ha5 == io_addra ? mem_165 : _GEN_164; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_166 = 8'ha6 == io_addra ? mem_166 : _GEN_165; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_167 = 8'ha7 == io_addra ? mem_167 : _GEN_166; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_168 = 8'ha8 == io_addra ? mem_168 : _GEN_167; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_169 = 8'ha9 == io_addra ? mem_169 : _GEN_168; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_170 = 8'haa == io_addra ? mem_170 : _GEN_169; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_171 = 8'hab == io_addra ? mem_171 : _GEN_170; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_172 = 8'hac == io_addra ? mem_172 : _GEN_171; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_173 = 8'had == io_addra ? mem_173 : _GEN_172; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_174 = 8'hae == io_addra ? mem_174 : _GEN_173; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_175 = 8'haf == io_addra ? mem_175 : _GEN_174; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_176 = 8'hb0 == io_addra ? mem_176 : _GEN_175; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_177 = 8'hb1 == io_addra ? mem_177 : _GEN_176; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_178 = 8'hb2 == io_addra ? mem_178 : _GEN_177; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_179 = 8'hb3 == io_addra ? mem_179 : _GEN_178; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_180 = 8'hb4 == io_addra ? mem_180 : _GEN_179; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_181 = 8'hb5 == io_addra ? mem_181 : _GEN_180; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_182 = 8'hb6 == io_addra ? mem_182 : _GEN_181; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_183 = 8'hb7 == io_addra ? mem_183 : _GEN_182; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_184 = 8'hb8 == io_addra ? mem_184 : _GEN_183; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_185 = 8'hb9 == io_addra ? mem_185 : _GEN_184; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_186 = 8'hba == io_addra ? mem_186 : _GEN_185; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_187 = 8'hbb == io_addra ? mem_187 : _GEN_186; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_188 = 8'hbc == io_addra ? mem_188 : _GEN_187; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_189 = 8'hbd == io_addra ? mem_189 : _GEN_188; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_190 = 8'hbe == io_addra ? mem_190 : _GEN_189; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_191 = 8'hbf == io_addra ? mem_191 : _GEN_190; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_192 = 8'hc0 == io_addra ? mem_192 : _GEN_191; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_193 = 8'hc1 == io_addra ? mem_193 : _GEN_192; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_194 = 8'hc2 == io_addra ? mem_194 : _GEN_193; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_195 = 8'hc3 == io_addra ? mem_195 : _GEN_194; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_196 = 8'hc4 == io_addra ? mem_196 : _GEN_195; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_197 = 8'hc5 == io_addra ? mem_197 : _GEN_196; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_198 = 8'hc6 == io_addra ? mem_198 : _GEN_197; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_199 = 8'hc7 == io_addra ? mem_199 : _GEN_198; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_200 = 8'hc8 == io_addra ? mem_200 : _GEN_199; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_201 = 8'hc9 == io_addra ? mem_201 : _GEN_200; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_202 = 8'hca == io_addra ? mem_202 : _GEN_201; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_203 = 8'hcb == io_addra ? mem_203 : _GEN_202; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_204 = 8'hcc == io_addra ? mem_204 : _GEN_203; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_205 = 8'hcd == io_addra ? mem_205 : _GEN_204; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_206 = 8'hce == io_addra ? mem_206 : _GEN_205; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_207 = 8'hcf == io_addra ? mem_207 : _GEN_206; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_208 = 8'hd0 == io_addra ? mem_208 : _GEN_207; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_209 = 8'hd1 == io_addra ? mem_209 : _GEN_208; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_210 = 8'hd2 == io_addra ? mem_210 : _GEN_209; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_211 = 8'hd3 == io_addra ? mem_211 : _GEN_210; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_212 = 8'hd4 == io_addra ? mem_212 : _GEN_211; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_213 = 8'hd5 == io_addra ? mem_213 : _GEN_212; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_214 = 8'hd6 == io_addra ? mem_214 : _GEN_213; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_215 = 8'hd7 == io_addra ? mem_215 : _GEN_214; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_216 = 8'hd8 == io_addra ? mem_216 : _GEN_215; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_217 = 8'hd9 == io_addra ? mem_217 : _GEN_216; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_218 = 8'hda == io_addra ? mem_218 : _GEN_217; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_219 = 8'hdb == io_addra ? mem_219 : _GEN_218; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_220 = 8'hdc == io_addra ? mem_220 : _GEN_219; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_221 = 8'hdd == io_addra ? mem_221 : _GEN_220; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_222 = 8'hde == io_addra ? mem_222 : _GEN_221; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_223 = 8'hdf == io_addra ? mem_223 : _GEN_222; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_224 = 8'he0 == io_addra ? mem_224 : _GEN_223; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_225 = 8'he1 == io_addra ? mem_225 : _GEN_224; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_226 = 8'he2 == io_addra ? mem_226 : _GEN_225; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_227 = 8'he3 == io_addra ? mem_227 : _GEN_226; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_228 = 8'he4 == io_addra ? mem_228 : _GEN_227; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_229 = 8'he5 == io_addra ? mem_229 : _GEN_228; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_230 = 8'he6 == io_addra ? mem_230 : _GEN_229; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_231 = 8'he7 == io_addra ? mem_231 : _GEN_230; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_232 = 8'he8 == io_addra ? mem_232 : _GEN_231; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_233 = 8'he9 == io_addra ? mem_233 : _GEN_232; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_234 = 8'hea == io_addra ? mem_234 : _GEN_233; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_235 = 8'heb == io_addra ? mem_235 : _GEN_234; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_236 = 8'hec == io_addra ? mem_236 : _GEN_235; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_237 = 8'hed == io_addra ? mem_237 : _GEN_236; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_238 = 8'hee == io_addra ? mem_238 : _GEN_237; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_239 = 8'hef == io_addra ? mem_239 : _GEN_238; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_240 = 8'hf0 == io_addra ? mem_240 : _GEN_239; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_241 = 8'hf1 == io_addra ? mem_241 : _GEN_240; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_242 = 8'hf2 == io_addra ? mem_242 : _GEN_241; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_243 = 8'hf3 == io_addra ? mem_243 : _GEN_242; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_244 = 8'hf4 == io_addra ? mem_244 : _GEN_243; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_245 = 8'hf5 == io_addra ? mem_245 : _GEN_244; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_246 = 8'hf6 == io_addra ? mem_246 : _GEN_245; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_247 = 8'hf7 == io_addra ? mem_247 : _GEN_246; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_248 = 8'hf8 == io_addra ? mem_248 : _GEN_247; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_249 = 8'hf9 == io_addra ? mem_249 : _GEN_248; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_250 = 8'hfa == io_addra ? mem_250 : _GEN_249; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [127:0] _GEN_251 = 8'hfb == io_addra ? mem_251 : _GEN_250; // @[RAM.scala 43:24 RAM.scala 43:24]
  assign io_douta = io_douta_REG; // @[RAM.scala 43:14]
  always @(posedge clock) begin
    if (reset) begin // @[RAM.scala 41:22]
      mem_0 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h0 == io_addrb) begin // @[RAM.scala 50:23]
        mem_0 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_1 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h1 == io_addrb) begin // @[RAM.scala 50:23]
        mem_1 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_2 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h2 == io_addrb) begin // @[RAM.scala 50:23]
        mem_2 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_3 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h3 == io_addrb) begin // @[RAM.scala 50:23]
        mem_3 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_4 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h4 == io_addrb) begin // @[RAM.scala 50:23]
        mem_4 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_5 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h5 == io_addrb) begin // @[RAM.scala 50:23]
        mem_5 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_6 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h6 == io_addrb) begin // @[RAM.scala 50:23]
        mem_6 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_7 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h7 == io_addrb) begin // @[RAM.scala 50:23]
        mem_7 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_8 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h8 == io_addrb) begin // @[RAM.scala 50:23]
        mem_8 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_9 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h9 == io_addrb) begin // @[RAM.scala 50:23]
        mem_9 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_10 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha == io_addrb) begin // @[RAM.scala 50:23]
        mem_10 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_11 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb == io_addrb) begin // @[RAM.scala 50:23]
        mem_11 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_12 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc == io_addrb) begin // @[RAM.scala 50:23]
        mem_12 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_13 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd == io_addrb) begin // @[RAM.scala 50:23]
        mem_13 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_14 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he == io_addrb) begin // @[RAM.scala 50:23]
        mem_14 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_15 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf == io_addrb) begin // @[RAM.scala 50:23]
        mem_15 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_16 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h10 == io_addrb) begin // @[RAM.scala 50:23]
        mem_16 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_17 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h11 == io_addrb) begin // @[RAM.scala 50:23]
        mem_17 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_18 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h12 == io_addrb) begin // @[RAM.scala 50:23]
        mem_18 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_19 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h13 == io_addrb) begin // @[RAM.scala 50:23]
        mem_19 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_20 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h14 == io_addrb) begin // @[RAM.scala 50:23]
        mem_20 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_21 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h15 == io_addrb) begin // @[RAM.scala 50:23]
        mem_21 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_22 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h16 == io_addrb) begin // @[RAM.scala 50:23]
        mem_22 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_23 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h17 == io_addrb) begin // @[RAM.scala 50:23]
        mem_23 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_24 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h18 == io_addrb) begin // @[RAM.scala 50:23]
        mem_24 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_25 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h19 == io_addrb) begin // @[RAM.scala 50:23]
        mem_25 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_26 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h1a == io_addrb) begin // @[RAM.scala 50:23]
        mem_26 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_27 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h1b == io_addrb) begin // @[RAM.scala 50:23]
        mem_27 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_28 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h1c == io_addrb) begin // @[RAM.scala 50:23]
        mem_28 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_29 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h1d == io_addrb) begin // @[RAM.scala 50:23]
        mem_29 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_30 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h1e == io_addrb) begin // @[RAM.scala 50:23]
        mem_30 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_31 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h1f == io_addrb) begin // @[RAM.scala 50:23]
        mem_31 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_32 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h20 == io_addrb) begin // @[RAM.scala 50:23]
        mem_32 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_33 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h21 == io_addrb) begin // @[RAM.scala 50:23]
        mem_33 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_34 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h22 == io_addrb) begin // @[RAM.scala 50:23]
        mem_34 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_35 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h23 == io_addrb) begin // @[RAM.scala 50:23]
        mem_35 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_36 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h24 == io_addrb) begin // @[RAM.scala 50:23]
        mem_36 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_37 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h25 == io_addrb) begin // @[RAM.scala 50:23]
        mem_37 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_38 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h26 == io_addrb) begin // @[RAM.scala 50:23]
        mem_38 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_39 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h27 == io_addrb) begin // @[RAM.scala 50:23]
        mem_39 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_40 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h28 == io_addrb) begin // @[RAM.scala 50:23]
        mem_40 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_41 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h29 == io_addrb) begin // @[RAM.scala 50:23]
        mem_41 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_42 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h2a == io_addrb) begin // @[RAM.scala 50:23]
        mem_42 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_43 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h2b == io_addrb) begin // @[RAM.scala 50:23]
        mem_43 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_44 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h2c == io_addrb) begin // @[RAM.scala 50:23]
        mem_44 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_45 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h2d == io_addrb) begin // @[RAM.scala 50:23]
        mem_45 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_46 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h2e == io_addrb) begin // @[RAM.scala 50:23]
        mem_46 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_47 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h2f == io_addrb) begin // @[RAM.scala 50:23]
        mem_47 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_48 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h30 == io_addrb) begin // @[RAM.scala 50:23]
        mem_48 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_49 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h31 == io_addrb) begin // @[RAM.scala 50:23]
        mem_49 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_50 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h32 == io_addrb) begin // @[RAM.scala 50:23]
        mem_50 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_51 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h33 == io_addrb) begin // @[RAM.scala 50:23]
        mem_51 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_52 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h34 == io_addrb) begin // @[RAM.scala 50:23]
        mem_52 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_53 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h35 == io_addrb) begin // @[RAM.scala 50:23]
        mem_53 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_54 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h36 == io_addrb) begin // @[RAM.scala 50:23]
        mem_54 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_55 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h37 == io_addrb) begin // @[RAM.scala 50:23]
        mem_55 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_56 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h38 == io_addrb) begin // @[RAM.scala 50:23]
        mem_56 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_57 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h39 == io_addrb) begin // @[RAM.scala 50:23]
        mem_57 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_58 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h3a == io_addrb) begin // @[RAM.scala 50:23]
        mem_58 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_59 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h3b == io_addrb) begin // @[RAM.scala 50:23]
        mem_59 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_60 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h3c == io_addrb) begin // @[RAM.scala 50:23]
        mem_60 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_61 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h3d == io_addrb) begin // @[RAM.scala 50:23]
        mem_61 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_62 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h3e == io_addrb) begin // @[RAM.scala 50:23]
        mem_62 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_63 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h3f == io_addrb) begin // @[RAM.scala 50:23]
        mem_63 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_64 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h40 == io_addrb) begin // @[RAM.scala 50:23]
        mem_64 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_65 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h41 == io_addrb) begin // @[RAM.scala 50:23]
        mem_65 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_66 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h42 == io_addrb) begin // @[RAM.scala 50:23]
        mem_66 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_67 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h43 == io_addrb) begin // @[RAM.scala 50:23]
        mem_67 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_68 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h44 == io_addrb) begin // @[RAM.scala 50:23]
        mem_68 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_69 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h45 == io_addrb) begin // @[RAM.scala 50:23]
        mem_69 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_70 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h46 == io_addrb) begin // @[RAM.scala 50:23]
        mem_70 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_71 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h47 == io_addrb) begin // @[RAM.scala 50:23]
        mem_71 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_72 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h48 == io_addrb) begin // @[RAM.scala 50:23]
        mem_72 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_73 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h49 == io_addrb) begin // @[RAM.scala 50:23]
        mem_73 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_74 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h4a == io_addrb) begin // @[RAM.scala 50:23]
        mem_74 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_75 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h4b == io_addrb) begin // @[RAM.scala 50:23]
        mem_75 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_76 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h4c == io_addrb) begin // @[RAM.scala 50:23]
        mem_76 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_77 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h4d == io_addrb) begin // @[RAM.scala 50:23]
        mem_77 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_78 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h4e == io_addrb) begin // @[RAM.scala 50:23]
        mem_78 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_79 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h4f == io_addrb) begin // @[RAM.scala 50:23]
        mem_79 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_80 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h50 == io_addrb) begin // @[RAM.scala 50:23]
        mem_80 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_81 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h51 == io_addrb) begin // @[RAM.scala 50:23]
        mem_81 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_82 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h52 == io_addrb) begin // @[RAM.scala 50:23]
        mem_82 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_83 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h53 == io_addrb) begin // @[RAM.scala 50:23]
        mem_83 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_84 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h54 == io_addrb) begin // @[RAM.scala 50:23]
        mem_84 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_85 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h55 == io_addrb) begin // @[RAM.scala 50:23]
        mem_85 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_86 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h56 == io_addrb) begin // @[RAM.scala 50:23]
        mem_86 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_87 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h57 == io_addrb) begin // @[RAM.scala 50:23]
        mem_87 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_88 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h58 == io_addrb) begin // @[RAM.scala 50:23]
        mem_88 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_89 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h59 == io_addrb) begin // @[RAM.scala 50:23]
        mem_89 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_90 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h5a == io_addrb) begin // @[RAM.scala 50:23]
        mem_90 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_91 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h5b == io_addrb) begin // @[RAM.scala 50:23]
        mem_91 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_92 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h5c == io_addrb) begin // @[RAM.scala 50:23]
        mem_92 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_93 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h5d == io_addrb) begin // @[RAM.scala 50:23]
        mem_93 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_94 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h5e == io_addrb) begin // @[RAM.scala 50:23]
        mem_94 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_95 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h5f == io_addrb) begin // @[RAM.scala 50:23]
        mem_95 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_96 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h60 == io_addrb) begin // @[RAM.scala 50:23]
        mem_96 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_97 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h61 == io_addrb) begin // @[RAM.scala 50:23]
        mem_97 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_98 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h62 == io_addrb) begin // @[RAM.scala 50:23]
        mem_98 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_99 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h63 == io_addrb) begin // @[RAM.scala 50:23]
        mem_99 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_100 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h64 == io_addrb) begin // @[RAM.scala 50:23]
        mem_100 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_101 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h65 == io_addrb) begin // @[RAM.scala 50:23]
        mem_101 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_102 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h66 == io_addrb) begin // @[RAM.scala 50:23]
        mem_102 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_103 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h67 == io_addrb) begin // @[RAM.scala 50:23]
        mem_103 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_104 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h68 == io_addrb) begin // @[RAM.scala 50:23]
        mem_104 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_105 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h69 == io_addrb) begin // @[RAM.scala 50:23]
        mem_105 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_106 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h6a == io_addrb) begin // @[RAM.scala 50:23]
        mem_106 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_107 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h6b == io_addrb) begin // @[RAM.scala 50:23]
        mem_107 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_108 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h6c == io_addrb) begin // @[RAM.scala 50:23]
        mem_108 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_109 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h6d == io_addrb) begin // @[RAM.scala 50:23]
        mem_109 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_110 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h6e == io_addrb) begin // @[RAM.scala 50:23]
        mem_110 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_111 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h6f == io_addrb) begin // @[RAM.scala 50:23]
        mem_111 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_112 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h70 == io_addrb) begin // @[RAM.scala 50:23]
        mem_112 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_113 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h71 == io_addrb) begin // @[RAM.scala 50:23]
        mem_113 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_114 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h72 == io_addrb) begin // @[RAM.scala 50:23]
        mem_114 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_115 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h73 == io_addrb) begin // @[RAM.scala 50:23]
        mem_115 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_116 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h74 == io_addrb) begin // @[RAM.scala 50:23]
        mem_116 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_117 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h75 == io_addrb) begin // @[RAM.scala 50:23]
        mem_117 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_118 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h76 == io_addrb) begin // @[RAM.scala 50:23]
        mem_118 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_119 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h77 == io_addrb) begin // @[RAM.scala 50:23]
        mem_119 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_120 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h78 == io_addrb) begin // @[RAM.scala 50:23]
        mem_120 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_121 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h79 == io_addrb) begin // @[RAM.scala 50:23]
        mem_121 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_122 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h7a == io_addrb) begin // @[RAM.scala 50:23]
        mem_122 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_123 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h7b == io_addrb) begin // @[RAM.scala 50:23]
        mem_123 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_124 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h7c == io_addrb) begin // @[RAM.scala 50:23]
        mem_124 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_125 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h7d == io_addrb) begin // @[RAM.scala 50:23]
        mem_125 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_126 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h7e == io_addrb) begin // @[RAM.scala 50:23]
        mem_126 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_127 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h7f == io_addrb) begin // @[RAM.scala 50:23]
        mem_127 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_128 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h80 == io_addrb) begin // @[RAM.scala 50:23]
        mem_128 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_129 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h81 == io_addrb) begin // @[RAM.scala 50:23]
        mem_129 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_130 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h82 == io_addrb) begin // @[RAM.scala 50:23]
        mem_130 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_131 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h83 == io_addrb) begin // @[RAM.scala 50:23]
        mem_131 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_132 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h84 == io_addrb) begin // @[RAM.scala 50:23]
        mem_132 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_133 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h85 == io_addrb) begin // @[RAM.scala 50:23]
        mem_133 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_134 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h86 == io_addrb) begin // @[RAM.scala 50:23]
        mem_134 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_135 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h87 == io_addrb) begin // @[RAM.scala 50:23]
        mem_135 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_136 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h88 == io_addrb) begin // @[RAM.scala 50:23]
        mem_136 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_137 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h89 == io_addrb) begin // @[RAM.scala 50:23]
        mem_137 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_138 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h8a == io_addrb) begin // @[RAM.scala 50:23]
        mem_138 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_139 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h8b == io_addrb) begin // @[RAM.scala 50:23]
        mem_139 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_140 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h8c == io_addrb) begin // @[RAM.scala 50:23]
        mem_140 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_141 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h8d == io_addrb) begin // @[RAM.scala 50:23]
        mem_141 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_142 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h8e == io_addrb) begin // @[RAM.scala 50:23]
        mem_142 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_143 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h8f == io_addrb) begin // @[RAM.scala 50:23]
        mem_143 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_144 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h90 == io_addrb) begin // @[RAM.scala 50:23]
        mem_144 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_145 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h91 == io_addrb) begin // @[RAM.scala 50:23]
        mem_145 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_146 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h92 == io_addrb) begin // @[RAM.scala 50:23]
        mem_146 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_147 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h93 == io_addrb) begin // @[RAM.scala 50:23]
        mem_147 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_148 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h94 == io_addrb) begin // @[RAM.scala 50:23]
        mem_148 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_149 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h95 == io_addrb) begin // @[RAM.scala 50:23]
        mem_149 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_150 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h96 == io_addrb) begin // @[RAM.scala 50:23]
        mem_150 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_151 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h97 == io_addrb) begin // @[RAM.scala 50:23]
        mem_151 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_152 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h98 == io_addrb) begin // @[RAM.scala 50:23]
        mem_152 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_153 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h99 == io_addrb) begin // @[RAM.scala 50:23]
        mem_153 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_154 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h9a == io_addrb) begin // @[RAM.scala 50:23]
        mem_154 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_155 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h9b == io_addrb) begin // @[RAM.scala 50:23]
        mem_155 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_156 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h9c == io_addrb) begin // @[RAM.scala 50:23]
        mem_156 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_157 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h9d == io_addrb) begin // @[RAM.scala 50:23]
        mem_157 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_158 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h9e == io_addrb) begin // @[RAM.scala 50:23]
        mem_158 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_159 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h9f == io_addrb) begin // @[RAM.scala 50:23]
        mem_159 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_160 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha0 == io_addrb) begin // @[RAM.scala 50:23]
        mem_160 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_161 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha1 == io_addrb) begin // @[RAM.scala 50:23]
        mem_161 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_162 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha2 == io_addrb) begin // @[RAM.scala 50:23]
        mem_162 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_163 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha3 == io_addrb) begin // @[RAM.scala 50:23]
        mem_163 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_164 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha4 == io_addrb) begin // @[RAM.scala 50:23]
        mem_164 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_165 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha5 == io_addrb) begin // @[RAM.scala 50:23]
        mem_165 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_166 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha6 == io_addrb) begin // @[RAM.scala 50:23]
        mem_166 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_167 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha7 == io_addrb) begin // @[RAM.scala 50:23]
        mem_167 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_168 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha8 == io_addrb) begin // @[RAM.scala 50:23]
        mem_168 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_169 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha9 == io_addrb) begin // @[RAM.scala 50:23]
        mem_169 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_170 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'haa == io_addrb) begin // @[RAM.scala 50:23]
        mem_170 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_171 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hab == io_addrb) begin // @[RAM.scala 50:23]
        mem_171 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_172 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hac == io_addrb) begin // @[RAM.scala 50:23]
        mem_172 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_173 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'had == io_addrb) begin // @[RAM.scala 50:23]
        mem_173 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_174 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hae == io_addrb) begin // @[RAM.scala 50:23]
        mem_174 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_175 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'haf == io_addrb) begin // @[RAM.scala 50:23]
        mem_175 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_176 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb0 == io_addrb) begin // @[RAM.scala 50:23]
        mem_176 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_177 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb1 == io_addrb) begin // @[RAM.scala 50:23]
        mem_177 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_178 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb2 == io_addrb) begin // @[RAM.scala 50:23]
        mem_178 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_179 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb3 == io_addrb) begin // @[RAM.scala 50:23]
        mem_179 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_180 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb4 == io_addrb) begin // @[RAM.scala 50:23]
        mem_180 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_181 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb5 == io_addrb) begin // @[RAM.scala 50:23]
        mem_181 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_182 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb6 == io_addrb) begin // @[RAM.scala 50:23]
        mem_182 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_183 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb7 == io_addrb) begin // @[RAM.scala 50:23]
        mem_183 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_184 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb8 == io_addrb) begin // @[RAM.scala 50:23]
        mem_184 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_185 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb9 == io_addrb) begin // @[RAM.scala 50:23]
        mem_185 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_186 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hba == io_addrb) begin // @[RAM.scala 50:23]
        mem_186 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_187 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hbb == io_addrb) begin // @[RAM.scala 50:23]
        mem_187 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_188 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hbc == io_addrb) begin // @[RAM.scala 50:23]
        mem_188 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_189 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hbd == io_addrb) begin // @[RAM.scala 50:23]
        mem_189 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_190 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hbe == io_addrb) begin // @[RAM.scala 50:23]
        mem_190 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_191 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hbf == io_addrb) begin // @[RAM.scala 50:23]
        mem_191 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_192 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc0 == io_addrb) begin // @[RAM.scala 50:23]
        mem_192 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_193 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc1 == io_addrb) begin // @[RAM.scala 50:23]
        mem_193 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_194 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc2 == io_addrb) begin // @[RAM.scala 50:23]
        mem_194 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_195 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc3 == io_addrb) begin // @[RAM.scala 50:23]
        mem_195 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_196 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc4 == io_addrb) begin // @[RAM.scala 50:23]
        mem_196 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_197 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc5 == io_addrb) begin // @[RAM.scala 50:23]
        mem_197 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_198 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc6 == io_addrb) begin // @[RAM.scala 50:23]
        mem_198 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_199 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc7 == io_addrb) begin // @[RAM.scala 50:23]
        mem_199 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_200 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc8 == io_addrb) begin // @[RAM.scala 50:23]
        mem_200 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_201 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc9 == io_addrb) begin // @[RAM.scala 50:23]
        mem_201 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_202 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hca == io_addrb) begin // @[RAM.scala 50:23]
        mem_202 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_203 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hcb == io_addrb) begin // @[RAM.scala 50:23]
        mem_203 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_204 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hcc == io_addrb) begin // @[RAM.scala 50:23]
        mem_204 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_205 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hcd == io_addrb) begin // @[RAM.scala 50:23]
        mem_205 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_206 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hce == io_addrb) begin // @[RAM.scala 50:23]
        mem_206 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_207 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hcf == io_addrb) begin // @[RAM.scala 50:23]
        mem_207 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_208 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd0 == io_addrb) begin // @[RAM.scala 50:23]
        mem_208 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_209 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd1 == io_addrb) begin // @[RAM.scala 50:23]
        mem_209 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_210 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd2 == io_addrb) begin // @[RAM.scala 50:23]
        mem_210 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_211 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd3 == io_addrb) begin // @[RAM.scala 50:23]
        mem_211 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_212 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd4 == io_addrb) begin // @[RAM.scala 50:23]
        mem_212 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_213 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd5 == io_addrb) begin // @[RAM.scala 50:23]
        mem_213 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_214 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd6 == io_addrb) begin // @[RAM.scala 50:23]
        mem_214 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_215 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd7 == io_addrb) begin // @[RAM.scala 50:23]
        mem_215 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_216 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd8 == io_addrb) begin // @[RAM.scala 50:23]
        mem_216 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_217 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd9 == io_addrb) begin // @[RAM.scala 50:23]
        mem_217 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_218 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hda == io_addrb) begin // @[RAM.scala 50:23]
        mem_218 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_219 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hdb == io_addrb) begin // @[RAM.scala 50:23]
        mem_219 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_220 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hdc == io_addrb) begin // @[RAM.scala 50:23]
        mem_220 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_221 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hdd == io_addrb) begin // @[RAM.scala 50:23]
        mem_221 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_222 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hde == io_addrb) begin // @[RAM.scala 50:23]
        mem_222 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_223 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hdf == io_addrb) begin // @[RAM.scala 50:23]
        mem_223 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_224 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he0 == io_addrb) begin // @[RAM.scala 50:23]
        mem_224 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_225 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he1 == io_addrb) begin // @[RAM.scala 50:23]
        mem_225 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_226 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he2 == io_addrb) begin // @[RAM.scala 50:23]
        mem_226 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_227 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he3 == io_addrb) begin // @[RAM.scala 50:23]
        mem_227 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_228 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he4 == io_addrb) begin // @[RAM.scala 50:23]
        mem_228 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_229 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he5 == io_addrb) begin // @[RAM.scala 50:23]
        mem_229 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_230 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he6 == io_addrb) begin // @[RAM.scala 50:23]
        mem_230 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_231 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he7 == io_addrb) begin // @[RAM.scala 50:23]
        mem_231 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_232 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he8 == io_addrb) begin // @[RAM.scala 50:23]
        mem_232 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_233 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he9 == io_addrb) begin // @[RAM.scala 50:23]
        mem_233 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_234 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hea == io_addrb) begin // @[RAM.scala 50:23]
        mem_234 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_235 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'heb == io_addrb) begin // @[RAM.scala 50:23]
        mem_235 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_236 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hec == io_addrb) begin // @[RAM.scala 50:23]
        mem_236 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_237 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hed == io_addrb) begin // @[RAM.scala 50:23]
        mem_237 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_238 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hee == io_addrb) begin // @[RAM.scala 50:23]
        mem_238 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_239 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hef == io_addrb) begin // @[RAM.scala 50:23]
        mem_239 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_240 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf0 == io_addrb) begin // @[RAM.scala 50:23]
        mem_240 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_241 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf1 == io_addrb) begin // @[RAM.scala 50:23]
        mem_241 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_242 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf2 == io_addrb) begin // @[RAM.scala 50:23]
        mem_242 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_243 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf3 == io_addrb) begin // @[RAM.scala 50:23]
        mem_243 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_244 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf4 == io_addrb) begin // @[RAM.scala 50:23]
        mem_244 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_245 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf5 == io_addrb) begin // @[RAM.scala 50:23]
        mem_245 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_246 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf6 == io_addrb) begin // @[RAM.scala 50:23]
        mem_246 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_247 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf7 == io_addrb) begin // @[RAM.scala 50:23]
        mem_247 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_248 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf8 == io_addrb) begin // @[RAM.scala 50:23]
        mem_248 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_249 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf9 == io_addrb) begin // @[RAM.scala 50:23]
        mem_249 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_250 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hfa == io_addrb) begin // @[RAM.scala 50:23]
        mem_250 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_251 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hfb == io_addrb) begin // @[RAM.scala 50:23]
        mem_251 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_252 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hfc == io_addrb) begin // @[RAM.scala 50:23]
        mem_252 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_253 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hfd == io_addrb) begin // @[RAM.scala 50:23]
        mem_253 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_254 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hfe == io_addrb) begin // @[RAM.scala 50:23]
        mem_254 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_255 <= 128'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hff == io_addrb) begin // @[RAM.scala 50:23]
        mem_255 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (8'hff == io_addra) begin // @[RAM.scala 43:24]
      io_douta_REG <= mem_255; // @[RAM.scala 43:24]
    end else if (8'hfe == io_addra) begin // @[RAM.scala 43:24]
      io_douta_REG <= mem_254; // @[RAM.scala 43:24]
    end else if (8'hfd == io_addra) begin // @[RAM.scala 43:24]
      io_douta_REG <= mem_253; // @[RAM.scala 43:24]
    end else if (8'hfc == io_addra) begin // @[RAM.scala 43:24]
      io_douta_REG <= mem_252; // @[RAM.scala 43:24]
    end else begin
      io_douta_REG <= _GEN_251;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  mem_0 = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  mem_1 = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  mem_2 = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  mem_3 = _RAND_3[127:0];
  _RAND_4 = {4{`RANDOM}};
  mem_4 = _RAND_4[127:0];
  _RAND_5 = {4{`RANDOM}};
  mem_5 = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  mem_6 = _RAND_6[127:0];
  _RAND_7 = {4{`RANDOM}};
  mem_7 = _RAND_7[127:0];
  _RAND_8 = {4{`RANDOM}};
  mem_8 = _RAND_8[127:0];
  _RAND_9 = {4{`RANDOM}};
  mem_9 = _RAND_9[127:0];
  _RAND_10 = {4{`RANDOM}};
  mem_10 = _RAND_10[127:0];
  _RAND_11 = {4{`RANDOM}};
  mem_11 = _RAND_11[127:0];
  _RAND_12 = {4{`RANDOM}};
  mem_12 = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  mem_13 = _RAND_13[127:0];
  _RAND_14 = {4{`RANDOM}};
  mem_14 = _RAND_14[127:0];
  _RAND_15 = {4{`RANDOM}};
  mem_15 = _RAND_15[127:0];
  _RAND_16 = {4{`RANDOM}};
  mem_16 = _RAND_16[127:0];
  _RAND_17 = {4{`RANDOM}};
  mem_17 = _RAND_17[127:0];
  _RAND_18 = {4{`RANDOM}};
  mem_18 = _RAND_18[127:0];
  _RAND_19 = {4{`RANDOM}};
  mem_19 = _RAND_19[127:0];
  _RAND_20 = {4{`RANDOM}};
  mem_20 = _RAND_20[127:0];
  _RAND_21 = {4{`RANDOM}};
  mem_21 = _RAND_21[127:0];
  _RAND_22 = {4{`RANDOM}};
  mem_22 = _RAND_22[127:0];
  _RAND_23 = {4{`RANDOM}};
  mem_23 = _RAND_23[127:0];
  _RAND_24 = {4{`RANDOM}};
  mem_24 = _RAND_24[127:0];
  _RAND_25 = {4{`RANDOM}};
  mem_25 = _RAND_25[127:0];
  _RAND_26 = {4{`RANDOM}};
  mem_26 = _RAND_26[127:0];
  _RAND_27 = {4{`RANDOM}};
  mem_27 = _RAND_27[127:0];
  _RAND_28 = {4{`RANDOM}};
  mem_28 = _RAND_28[127:0];
  _RAND_29 = {4{`RANDOM}};
  mem_29 = _RAND_29[127:0];
  _RAND_30 = {4{`RANDOM}};
  mem_30 = _RAND_30[127:0];
  _RAND_31 = {4{`RANDOM}};
  mem_31 = _RAND_31[127:0];
  _RAND_32 = {4{`RANDOM}};
  mem_32 = _RAND_32[127:0];
  _RAND_33 = {4{`RANDOM}};
  mem_33 = _RAND_33[127:0];
  _RAND_34 = {4{`RANDOM}};
  mem_34 = _RAND_34[127:0];
  _RAND_35 = {4{`RANDOM}};
  mem_35 = _RAND_35[127:0];
  _RAND_36 = {4{`RANDOM}};
  mem_36 = _RAND_36[127:0];
  _RAND_37 = {4{`RANDOM}};
  mem_37 = _RAND_37[127:0];
  _RAND_38 = {4{`RANDOM}};
  mem_38 = _RAND_38[127:0];
  _RAND_39 = {4{`RANDOM}};
  mem_39 = _RAND_39[127:0];
  _RAND_40 = {4{`RANDOM}};
  mem_40 = _RAND_40[127:0];
  _RAND_41 = {4{`RANDOM}};
  mem_41 = _RAND_41[127:0];
  _RAND_42 = {4{`RANDOM}};
  mem_42 = _RAND_42[127:0];
  _RAND_43 = {4{`RANDOM}};
  mem_43 = _RAND_43[127:0];
  _RAND_44 = {4{`RANDOM}};
  mem_44 = _RAND_44[127:0];
  _RAND_45 = {4{`RANDOM}};
  mem_45 = _RAND_45[127:0];
  _RAND_46 = {4{`RANDOM}};
  mem_46 = _RAND_46[127:0];
  _RAND_47 = {4{`RANDOM}};
  mem_47 = _RAND_47[127:0];
  _RAND_48 = {4{`RANDOM}};
  mem_48 = _RAND_48[127:0];
  _RAND_49 = {4{`RANDOM}};
  mem_49 = _RAND_49[127:0];
  _RAND_50 = {4{`RANDOM}};
  mem_50 = _RAND_50[127:0];
  _RAND_51 = {4{`RANDOM}};
  mem_51 = _RAND_51[127:0];
  _RAND_52 = {4{`RANDOM}};
  mem_52 = _RAND_52[127:0];
  _RAND_53 = {4{`RANDOM}};
  mem_53 = _RAND_53[127:0];
  _RAND_54 = {4{`RANDOM}};
  mem_54 = _RAND_54[127:0];
  _RAND_55 = {4{`RANDOM}};
  mem_55 = _RAND_55[127:0];
  _RAND_56 = {4{`RANDOM}};
  mem_56 = _RAND_56[127:0];
  _RAND_57 = {4{`RANDOM}};
  mem_57 = _RAND_57[127:0];
  _RAND_58 = {4{`RANDOM}};
  mem_58 = _RAND_58[127:0];
  _RAND_59 = {4{`RANDOM}};
  mem_59 = _RAND_59[127:0];
  _RAND_60 = {4{`RANDOM}};
  mem_60 = _RAND_60[127:0];
  _RAND_61 = {4{`RANDOM}};
  mem_61 = _RAND_61[127:0];
  _RAND_62 = {4{`RANDOM}};
  mem_62 = _RAND_62[127:0];
  _RAND_63 = {4{`RANDOM}};
  mem_63 = _RAND_63[127:0];
  _RAND_64 = {4{`RANDOM}};
  mem_64 = _RAND_64[127:0];
  _RAND_65 = {4{`RANDOM}};
  mem_65 = _RAND_65[127:0];
  _RAND_66 = {4{`RANDOM}};
  mem_66 = _RAND_66[127:0];
  _RAND_67 = {4{`RANDOM}};
  mem_67 = _RAND_67[127:0];
  _RAND_68 = {4{`RANDOM}};
  mem_68 = _RAND_68[127:0];
  _RAND_69 = {4{`RANDOM}};
  mem_69 = _RAND_69[127:0];
  _RAND_70 = {4{`RANDOM}};
  mem_70 = _RAND_70[127:0];
  _RAND_71 = {4{`RANDOM}};
  mem_71 = _RAND_71[127:0];
  _RAND_72 = {4{`RANDOM}};
  mem_72 = _RAND_72[127:0];
  _RAND_73 = {4{`RANDOM}};
  mem_73 = _RAND_73[127:0];
  _RAND_74 = {4{`RANDOM}};
  mem_74 = _RAND_74[127:0];
  _RAND_75 = {4{`RANDOM}};
  mem_75 = _RAND_75[127:0];
  _RAND_76 = {4{`RANDOM}};
  mem_76 = _RAND_76[127:0];
  _RAND_77 = {4{`RANDOM}};
  mem_77 = _RAND_77[127:0];
  _RAND_78 = {4{`RANDOM}};
  mem_78 = _RAND_78[127:0];
  _RAND_79 = {4{`RANDOM}};
  mem_79 = _RAND_79[127:0];
  _RAND_80 = {4{`RANDOM}};
  mem_80 = _RAND_80[127:0];
  _RAND_81 = {4{`RANDOM}};
  mem_81 = _RAND_81[127:0];
  _RAND_82 = {4{`RANDOM}};
  mem_82 = _RAND_82[127:0];
  _RAND_83 = {4{`RANDOM}};
  mem_83 = _RAND_83[127:0];
  _RAND_84 = {4{`RANDOM}};
  mem_84 = _RAND_84[127:0];
  _RAND_85 = {4{`RANDOM}};
  mem_85 = _RAND_85[127:0];
  _RAND_86 = {4{`RANDOM}};
  mem_86 = _RAND_86[127:0];
  _RAND_87 = {4{`RANDOM}};
  mem_87 = _RAND_87[127:0];
  _RAND_88 = {4{`RANDOM}};
  mem_88 = _RAND_88[127:0];
  _RAND_89 = {4{`RANDOM}};
  mem_89 = _RAND_89[127:0];
  _RAND_90 = {4{`RANDOM}};
  mem_90 = _RAND_90[127:0];
  _RAND_91 = {4{`RANDOM}};
  mem_91 = _RAND_91[127:0];
  _RAND_92 = {4{`RANDOM}};
  mem_92 = _RAND_92[127:0];
  _RAND_93 = {4{`RANDOM}};
  mem_93 = _RAND_93[127:0];
  _RAND_94 = {4{`RANDOM}};
  mem_94 = _RAND_94[127:0];
  _RAND_95 = {4{`RANDOM}};
  mem_95 = _RAND_95[127:0];
  _RAND_96 = {4{`RANDOM}};
  mem_96 = _RAND_96[127:0];
  _RAND_97 = {4{`RANDOM}};
  mem_97 = _RAND_97[127:0];
  _RAND_98 = {4{`RANDOM}};
  mem_98 = _RAND_98[127:0];
  _RAND_99 = {4{`RANDOM}};
  mem_99 = _RAND_99[127:0];
  _RAND_100 = {4{`RANDOM}};
  mem_100 = _RAND_100[127:0];
  _RAND_101 = {4{`RANDOM}};
  mem_101 = _RAND_101[127:0];
  _RAND_102 = {4{`RANDOM}};
  mem_102 = _RAND_102[127:0];
  _RAND_103 = {4{`RANDOM}};
  mem_103 = _RAND_103[127:0];
  _RAND_104 = {4{`RANDOM}};
  mem_104 = _RAND_104[127:0];
  _RAND_105 = {4{`RANDOM}};
  mem_105 = _RAND_105[127:0];
  _RAND_106 = {4{`RANDOM}};
  mem_106 = _RAND_106[127:0];
  _RAND_107 = {4{`RANDOM}};
  mem_107 = _RAND_107[127:0];
  _RAND_108 = {4{`RANDOM}};
  mem_108 = _RAND_108[127:0];
  _RAND_109 = {4{`RANDOM}};
  mem_109 = _RAND_109[127:0];
  _RAND_110 = {4{`RANDOM}};
  mem_110 = _RAND_110[127:0];
  _RAND_111 = {4{`RANDOM}};
  mem_111 = _RAND_111[127:0];
  _RAND_112 = {4{`RANDOM}};
  mem_112 = _RAND_112[127:0];
  _RAND_113 = {4{`RANDOM}};
  mem_113 = _RAND_113[127:0];
  _RAND_114 = {4{`RANDOM}};
  mem_114 = _RAND_114[127:0];
  _RAND_115 = {4{`RANDOM}};
  mem_115 = _RAND_115[127:0];
  _RAND_116 = {4{`RANDOM}};
  mem_116 = _RAND_116[127:0];
  _RAND_117 = {4{`RANDOM}};
  mem_117 = _RAND_117[127:0];
  _RAND_118 = {4{`RANDOM}};
  mem_118 = _RAND_118[127:0];
  _RAND_119 = {4{`RANDOM}};
  mem_119 = _RAND_119[127:0];
  _RAND_120 = {4{`RANDOM}};
  mem_120 = _RAND_120[127:0];
  _RAND_121 = {4{`RANDOM}};
  mem_121 = _RAND_121[127:0];
  _RAND_122 = {4{`RANDOM}};
  mem_122 = _RAND_122[127:0];
  _RAND_123 = {4{`RANDOM}};
  mem_123 = _RAND_123[127:0];
  _RAND_124 = {4{`RANDOM}};
  mem_124 = _RAND_124[127:0];
  _RAND_125 = {4{`RANDOM}};
  mem_125 = _RAND_125[127:0];
  _RAND_126 = {4{`RANDOM}};
  mem_126 = _RAND_126[127:0];
  _RAND_127 = {4{`RANDOM}};
  mem_127 = _RAND_127[127:0];
  _RAND_128 = {4{`RANDOM}};
  mem_128 = _RAND_128[127:0];
  _RAND_129 = {4{`RANDOM}};
  mem_129 = _RAND_129[127:0];
  _RAND_130 = {4{`RANDOM}};
  mem_130 = _RAND_130[127:0];
  _RAND_131 = {4{`RANDOM}};
  mem_131 = _RAND_131[127:0];
  _RAND_132 = {4{`RANDOM}};
  mem_132 = _RAND_132[127:0];
  _RAND_133 = {4{`RANDOM}};
  mem_133 = _RAND_133[127:0];
  _RAND_134 = {4{`RANDOM}};
  mem_134 = _RAND_134[127:0];
  _RAND_135 = {4{`RANDOM}};
  mem_135 = _RAND_135[127:0];
  _RAND_136 = {4{`RANDOM}};
  mem_136 = _RAND_136[127:0];
  _RAND_137 = {4{`RANDOM}};
  mem_137 = _RAND_137[127:0];
  _RAND_138 = {4{`RANDOM}};
  mem_138 = _RAND_138[127:0];
  _RAND_139 = {4{`RANDOM}};
  mem_139 = _RAND_139[127:0];
  _RAND_140 = {4{`RANDOM}};
  mem_140 = _RAND_140[127:0];
  _RAND_141 = {4{`RANDOM}};
  mem_141 = _RAND_141[127:0];
  _RAND_142 = {4{`RANDOM}};
  mem_142 = _RAND_142[127:0];
  _RAND_143 = {4{`RANDOM}};
  mem_143 = _RAND_143[127:0];
  _RAND_144 = {4{`RANDOM}};
  mem_144 = _RAND_144[127:0];
  _RAND_145 = {4{`RANDOM}};
  mem_145 = _RAND_145[127:0];
  _RAND_146 = {4{`RANDOM}};
  mem_146 = _RAND_146[127:0];
  _RAND_147 = {4{`RANDOM}};
  mem_147 = _RAND_147[127:0];
  _RAND_148 = {4{`RANDOM}};
  mem_148 = _RAND_148[127:0];
  _RAND_149 = {4{`RANDOM}};
  mem_149 = _RAND_149[127:0];
  _RAND_150 = {4{`RANDOM}};
  mem_150 = _RAND_150[127:0];
  _RAND_151 = {4{`RANDOM}};
  mem_151 = _RAND_151[127:0];
  _RAND_152 = {4{`RANDOM}};
  mem_152 = _RAND_152[127:0];
  _RAND_153 = {4{`RANDOM}};
  mem_153 = _RAND_153[127:0];
  _RAND_154 = {4{`RANDOM}};
  mem_154 = _RAND_154[127:0];
  _RAND_155 = {4{`RANDOM}};
  mem_155 = _RAND_155[127:0];
  _RAND_156 = {4{`RANDOM}};
  mem_156 = _RAND_156[127:0];
  _RAND_157 = {4{`RANDOM}};
  mem_157 = _RAND_157[127:0];
  _RAND_158 = {4{`RANDOM}};
  mem_158 = _RAND_158[127:0];
  _RAND_159 = {4{`RANDOM}};
  mem_159 = _RAND_159[127:0];
  _RAND_160 = {4{`RANDOM}};
  mem_160 = _RAND_160[127:0];
  _RAND_161 = {4{`RANDOM}};
  mem_161 = _RAND_161[127:0];
  _RAND_162 = {4{`RANDOM}};
  mem_162 = _RAND_162[127:0];
  _RAND_163 = {4{`RANDOM}};
  mem_163 = _RAND_163[127:0];
  _RAND_164 = {4{`RANDOM}};
  mem_164 = _RAND_164[127:0];
  _RAND_165 = {4{`RANDOM}};
  mem_165 = _RAND_165[127:0];
  _RAND_166 = {4{`RANDOM}};
  mem_166 = _RAND_166[127:0];
  _RAND_167 = {4{`RANDOM}};
  mem_167 = _RAND_167[127:0];
  _RAND_168 = {4{`RANDOM}};
  mem_168 = _RAND_168[127:0];
  _RAND_169 = {4{`RANDOM}};
  mem_169 = _RAND_169[127:0];
  _RAND_170 = {4{`RANDOM}};
  mem_170 = _RAND_170[127:0];
  _RAND_171 = {4{`RANDOM}};
  mem_171 = _RAND_171[127:0];
  _RAND_172 = {4{`RANDOM}};
  mem_172 = _RAND_172[127:0];
  _RAND_173 = {4{`RANDOM}};
  mem_173 = _RAND_173[127:0];
  _RAND_174 = {4{`RANDOM}};
  mem_174 = _RAND_174[127:0];
  _RAND_175 = {4{`RANDOM}};
  mem_175 = _RAND_175[127:0];
  _RAND_176 = {4{`RANDOM}};
  mem_176 = _RAND_176[127:0];
  _RAND_177 = {4{`RANDOM}};
  mem_177 = _RAND_177[127:0];
  _RAND_178 = {4{`RANDOM}};
  mem_178 = _RAND_178[127:0];
  _RAND_179 = {4{`RANDOM}};
  mem_179 = _RAND_179[127:0];
  _RAND_180 = {4{`RANDOM}};
  mem_180 = _RAND_180[127:0];
  _RAND_181 = {4{`RANDOM}};
  mem_181 = _RAND_181[127:0];
  _RAND_182 = {4{`RANDOM}};
  mem_182 = _RAND_182[127:0];
  _RAND_183 = {4{`RANDOM}};
  mem_183 = _RAND_183[127:0];
  _RAND_184 = {4{`RANDOM}};
  mem_184 = _RAND_184[127:0];
  _RAND_185 = {4{`RANDOM}};
  mem_185 = _RAND_185[127:0];
  _RAND_186 = {4{`RANDOM}};
  mem_186 = _RAND_186[127:0];
  _RAND_187 = {4{`RANDOM}};
  mem_187 = _RAND_187[127:0];
  _RAND_188 = {4{`RANDOM}};
  mem_188 = _RAND_188[127:0];
  _RAND_189 = {4{`RANDOM}};
  mem_189 = _RAND_189[127:0];
  _RAND_190 = {4{`RANDOM}};
  mem_190 = _RAND_190[127:0];
  _RAND_191 = {4{`RANDOM}};
  mem_191 = _RAND_191[127:0];
  _RAND_192 = {4{`RANDOM}};
  mem_192 = _RAND_192[127:0];
  _RAND_193 = {4{`RANDOM}};
  mem_193 = _RAND_193[127:0];
  _RAND_194 = {4{`RANDOM}};
  mem_194 = _RAND_194[127:0];
  _RAND_195 = {4{`RANDOM}};
  mem_195 = _RAND_195[127:0];
  _RAND_196 = {4{`RANDOM}};
  mem_196 = _RAND_196[127:0];
  _RAND_197 = {4{`RANDOM}};
  mem_197 = _RAND_197[127:0];
  _RAND_198 = {4{`RANDOM}};
  mem_198 = _RAND_198[127:0];
  _RAND_199 = {4{`RANDOM}};
  mem_199 = _RAND_199[127:0];
  _RAND_200 = {4{`RANDOM}};
  mem_200 = _RAND_200[127:0];
  _RAND_201 = {4{`RANDOM}};
  mem_201 = _RAND_201[127:0];
  _RAND_202 = {4{`RANDOM}};
  mem_202 = _RAND_202[127:0];
  _RAND_203 = {4{`RANDOM}};
  mem_203 = _RAND_203[127:0];
  _RAND_204 = {4{`RANDOM}};
  mem_204 = _RAND_204[127:0];
  _RAND_205 = {4{`RANDOM}};
  mem_205 = _RAND_205[127:0];
  _RAND_206 = {4{`RANDOM}};
  mem_206 = _RAND_206[127:0];
  _RAND_207 = {4{`RANDOM}};
  mem_207 = _RAND_207[127:0];
  _RAND_208 = {4{`RANDOM}};
  mem_208 = _RAND_208[127:0];
  _RAND_209 = {4{`RANDOM}};
  mem_209 = _RAND_209[127:0];
  _RAND_210 = {4{`RANDOM}};
  mem_210 = _RAND_210[127:0];
  _RAND_211 = {4{`RANDOM}};
  mem_211 = _RAND_211[127:0];
  _RAND_212 = {4{`RANDOM}};
  mem_212 = _RAND_212[127:0];
  _RAND_213 = {4{`RANDOM}};
  mem_213 = _RAND_213[127:0];
  _RAND_214 = {4{`RANDOM}};
  mem_214 = _RAND_214[127:0];
  _RAND_215 = {4{`RANDOM}};
  mem_215 = _RAND_215[127:0];
  _RAND_216 = {4{`RANDOM}};
  mem_216 = _RAND_216[127:0];
  _RAND_217 = {4{`RANDOM}};
  mem_217 = _RAND_217[127:0];
  _RAND_218 = {4{`RANDOM}};
  mem_218 = _RAND_218[127:0];
  _RAND_219 = {4{`RANDOM}};
  mem_219 = _RAND_219[127:0];
  _RAND_220 = {4{`RANDOM}};
  mem_220 = _RAND_220[127:0];
  _RAND_221 = {4{`RANDOM}};
  mem_221 = _RAND_221[127:0];
  _RAND_222 = {4{`RANDOM}};
  mem_222 = _RAND_222[127:0];
  _RAND_223 = {4{`RANDOM}};
  mem_223 = _RAND_223[127:0];
  _RAND_224 = {4{`RANDOM}};
  mem_224 = _RAND_224[127:0];
  _RAND_225 = {4{`RANDOM}};
  mem_225 = _RAND_225[127:0];
  _RAND_226 = {4{`RANDOM}};
  mem_226 = _RAND_226[127:0];
  _RAND_227 = {4{`RANDOM}};
  mem_227 = _RAND_227[127:0];
  _RAND_228 = {4{`RANDOM}};
  mem_228 = _RAND_228[127:0];
  _RAND_229 = {4{`RANDOM}};
  mem_229 = _RAND_229[127:0];
  _RAND_230 = {4{`RANDOM}};
  mem_230 = _RAND_230[127:0];
  _RAND_231 = {4{`RANDOM}};
  mem_231 = _RAND_231[127:0];
  _RAND_232 = {4{`RANDOM}};
  mem_232 = _RAND_232[127:0];
  _RAND_233 = {4{`RANDOM}};
  mem_233 = _RAND_233[127:0];
  _RAND_234 = {4{`RANDOM}};
  mem_234 = _RAND_234[127:0];
  _RAND_235 = {4{`RANDOM}};
  mem_235 = _RAND_235[127:0];
  _RAND_236 = {4{`RANDOM}};
  mem_236 = _RAND_236[127:0];
  _RAND_237 = {4{`RANDOM}};
  mem_237 = _RAND_237[127:0];
  _RAND_238 = {4{`RANDOM}};
  mem_238 = _RAND_238[127:0];
  _RAND_239 = {4{`RANDOM}};
  mem_239 = _RAND_239[127:0];
  _RAND_240 = {4{`RANDOM}};
  mem_240 = _RAND_240[127:0];
  _RAND_241 = {4{`RANDOM}};
  mem_241 = _RAND_241[127:0];
  _RAND_242 = {4{`RANDOM}};
  mem_242 = _RAND_242[127:0];
  _RAND_243 = {4{`RANDOM}};
  mem_243 = _RAND_243[127:0];
  _RAND_244 = {4{`RANDOM}};
  mem_244 = _RAND_244[127:0];
  _RAND_245 = {4{`RANDOM}};
  mem_245 = _RAND_245[127:0];
  _RAND_246 = {4{`RANDOM}};
  mem_246 = _RAND_246[127:0];
  _RAND_247 = {4{`RANDOM}};
  mem_247 = _RAND_247[127:0];
  _RAND_248 = {4{`RANDOM}};
  mem_248 = _RAND_248[127:0];
  _RAND_249 = {4{`RANDOM}};
  mem_249 = _RAND_249[127:0];
  _RAND_250 = {4{`RANDOM}};
  mem_250 = _RAND_250[127:0];
  _RAND_251 = {4{`RANDOM}};
  mem_251 = _RAND_251[127:0];
  _RAND_252 = {4{`RANDOM}};
  mem_252 = _RAND_252[127:0];
  _RAND_253 = {4{`RANDOM}};
  mem_253 = _RAND_253[127:0];
  _RAND_254 = {4{`RANDOM}};
  mem_254 = _RAND_254[127:0];
  _RAND_255 = {4{`RANDOM}};
  mem_255 = _RAND_255[127:0];
  _RAND_256 = {4{`RANDOM}};
  io_douta_REG = _RAND_256[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DualPortBRAM(
  input          clock,
  input          reset,
  input          io_web,
  input  [7:0]   io_addra,
  input  [7:0]   io_addrb,
  input  [127:0] io_dinb,
  output [127:0] io_douta
);
  wire  sim_dual_port_bram_clock; // @[RAM.scala 30:40]
  wire  sim_dual_port_bram_reset; // @[RAM.scala 30:40]
  wire  sim_dual_port_bram_io_web; // @[RAM.scala 30:40]
  wire [7:0] sim_dual_port_bram_io_addra; // @[RAM.scala 30:40]
  wire [7:0] sim_dual_port_bram_io_addrb; // @[RAM.scala 30:40]
  wire [127:0] sim_dual_port_bram_io_dinb; // @[RAM.scala 30:40]
  wire [127:0] sim_dual_port_bram_io_douta; // @[RAM.scala 30:40]
  SimDualPortBRAM sim_dual_port_bram ( // @[RAM.scala 30:40]
    .clock(sim_dual_port_bram_clock),
    .reset(sim_dual_port_bram_reset),
    .io_web(sim_dual_port_bram_io_web),
    .io_addra(sim_dual_port_bram_io_addra),
    .io_addrb(sim_dual_port_bram_io_addrb),
    .io_dinb(sim_dual_port_bram_io_dinb),
    .io_douta(sim_dual_port_bram_io_douta)
  );
  assign io_douta = sim_dual_port_bram_io_douta; // @[RAM.scala 31:31]
  assign sim_dual_port_bram_clock = clock;
  assign sim_dual_port_bram_reset = reset;
  assign sim_dual_port_bram_io_web = io_web; // @[RAM.scala 31:31]
  assign sim_dual_port_bram_io_addra = io_addra; // @[RAM.scala 31:31]
  assign sim_dual_port_bram_io_addrb = io_addrb; // @[RAM.scala 31:31]
  assign sim_dual_port_bram_io_dinb = io_dinb; // @[RAM.scala 31:31]
endmodule
module SimDualPortBRAM_2(
  input         clock,
  input         reset,
  input         io_web,
  input  [7:0]  io_addra,
  input  [7:0]  io_addrb,
  input  [21:0] io_dinb,
  output [21:0] io_douta
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
`endif // RANDOMIZE_REG_INIT
  reg [21:0] mem_0; // @[RAM.scala 41:22]
  reg [21:0] mem_1; // @[RAM.scala 41:22]
  reg [21:0] mem_2; // @[RAM.scala 41:22]
  reg [21:0] mem_3; // @[RAM.scala 41:22]
  reg [21:0] mem_4; // @[RAM.scala 41:22]
  reg [21:0] mem_5; // @[RAM.scala 41:22]
  reg [21:0] mem_6; // @[RAM.scala 41:22]
  reg [21:0] mem_7; // @[RAM.scala 41:22]
  reg [21:0] mem_8; // @[RAM.scala 41:22]
  reg [21:0] mem_9; // @[RAM.scala 41:22]
  reg [21:0] mem_10; // @[RAM.scala 41:22]
  reg [21:0] mem_11; // @[RAM.scala 41:22]
  reg [21:0] mem_12; // @[RAM.scala 41:22]
  reg [21:0] mem_13; // @[RAM.scala 41:22]
  reg [21:0] mem_14; // @[RAM.scala 41:22]
  reg [21:0] mem_15; // @[RAM.scala 41:22]
  reg [21:0] mem_16; // @[RAM.scala 41:22]
  reg [21:0] mem_17; // @[RAM.scala 41:22]
  reg [21:0] mem_18; // @[RAM.scala 41:22]
  reg [21:0] mem_19; // @[RAM.scala 41:22]
  reg [21:0] mem_20; // @[RAM.scala 41:22]
  reg [21:0] mem_21; // @[RAM.scala 41:22]
  reg [21:0] mem_22; // @[RAM.scala 41:22]
  reg [21:0] mem_23; // @[RAM.scala 41:22]
  reg [21:0] mem_24; // @[RAM.scala 41:22]
  reg [21:0] mem_25; // @[RAM.scala 41:22]
  reg [21:0] mem_26; // @[RAM.scala 41:22]
  reg [21:0] mem_27; // @[RAM.scala 41:22]
  reg [21:0] mem_28; // @[RAM.scala 41:22]
  reg [21:0] mem_29; // @[RAM.scala 41:22]
  reg [21:0] mem_30; // @[RAM.scala 41:22]
  reg [21:0] mem_31; // @[RAM.scala 41:22]
  reg [21:0] mem_32; // @[RAM.scala 41:22]
  reg [21:0] mem_33; // @[RAM.scala 41:22]
  reg [21:0] mem_34; // @[RAM.scala 41:22]
  reg [21:0] mem_35; // @[RAM.scala 41:22]
  reg [21:0] mem_36; // @[RAM.scala 41:22]
  reg [21:0] mem_37; // @[RAM.scala 41:22]
  reg [21:0] mem_38; // @[RAM.scala 41:22]
  reg [21:0] mem_39; // @[RAM.scala 41:22]
  reg [21:0] mem_40; // @[RAM.scala 41:22]
  reg [21:0] mem_41; // @[RAM.scala 41:22]
  reg [21:0] mem_42; // @[RAM.scala 41:22]
  reg [21:0] mem_43; // @[RAM.scala 41:22]
  reg [21:0] mem_44; // @[RAM.scala 41:22]
  reg [21:0] mem_45; // @[RAM.scala 41:22]
  reg [21:0] mem_46; // @[RAM.scala 41:22]
  reg [21:0] mem_47; // @[RAM.scala 41:22]
  reg [21:0] mem_48; // @[RAM.scala 41:22]
  reg [21:0] mem_49; // @[RAM.scala 41:22]
  reg [21:0] mem_50; // @[RAM.scala 41:22]
  reg [21:0] mem_51; // @[RAM.scala 41:22]
  reg [21:0] mem_52; // @[RAM.scala 41:22]
  reg [21:0] mem_53; // @[RAM.scala 41:22]
  reg [21:0] mem_54; // @[RAM.scala 41:22]
  reg [21:0] mem_55; // @[RAM.scala 41:22]
  reg [21:0] mem_56; // @[RAM.scala 41:22]
  reg [21:0] mem_57; // @[RAM.scala 41:22]
  reg [21:0] mem_58; // @[RAM.scala 41:22]
  reg [21:0] mem_59; // @[RAM.scala 41:22]
  reg [21:0] mem_60; // @[RAM.scala 41:22]
  reg [21:0] mem_61; // @[RAM.scala 41:22]
  reg [21:0] mem_62; // @[RAM.scala 41:22]
  reg [21:0] mem_63; // @[RAM.scala 41:22]
  reg [21:0] mem_64; // @[RAM.scala 41:22]
  reg [21:0] mem_65; // @[RAM.scala 41:22]
  reg [21:0] mem_66; // @[RAM.scala 41:22]
  reg [21:0] mem_67; // @[RAM.scala 41:22]
  reg [21:0] mem_68; // @[RAM.scala 41:22]
  reg [21:0] mem_69; // @[RAM.scala 41:22]
  reg [21:0] mem_70; // @[RAM.scala 41:22]
  reg [21:0] mem_71; // @[RAM.scala 41:22]
  reg [21:0] mem_72; // @[RAM.scala 41:22]
  reg [21:0] mem_73; // @[RAM.scala 41:22]
  reg [21:0] mem_74; // @[RAM.scala 41:22]
  reg [21:0] mem_75; // @[RAM.scala 41:22]
  reg [21:0] mem_76; // @[RAM.scala 41:22]
  reg [21:0] mem_77; // @[RAM.scala 41:22]
  reg [21:0] mem_78; // @[RAM.scala 41:22]
  reg [21:0] mem_79; // @[RAM.scala 41:22]
  reg [21:0] mem_80; // @[RAM.scala 41:22]
  reg [21:0] mem_81; // @[RAM.scala 41:22]
  reg [21:0] mem_82; // @[RAM.scala 41:22]
  reg [21:0] mem_83; // @[RAM.scala 41:22]
  reg [21:0] mem_84; // @[RAM.scala 41:22]
  reg [21:0] mem_85; // @[RAM.scala 41:22]
  reg [21:0] mem_86; // @[RAM.scala 41:22]
  reg [21:0] mem_87; // @[RAM.scala 41:22]
  reg [21:0] mem_88; // @[RAM.scala 41:22]
  reg [21:0] mem_89; // @[RAM.scala 41:22]
  reg [21:0] mem_90; // @[RAM.scala 41:22]
  reg [21:0] mem_91; // @[RAM.scala 41:22]
  reg [21:0] mem_92; // @[RAM.scala 41:22]
  reg [21:0] mem_93; // @[RAM.scala 41:22]
  reg [21:0] mem_94; // @[RAM.scala 41:22]
  reg [21:0] mem_95; // @[RAM.scala 41:22]
  reg [21:0] mem_96; // @[RAM.scala 41:22]
  reg [21:0] mem_97; // @[RAM.scala 41:22]
  reg [21:0] mem_98; // @[RAM.scala 41:22]
  reg [21:0] mem_99; // @[RAM.scala 41:22]
  reg [21:0] mem_100; // @[RAM.scala 41:22]
  reg [21:0] mem_101; // @[RAM.scala 41:22]
  reg [21:0] mem_102; // @[RAM.scala 41:22]
  reg [21:0] mem_103; // @[RAM.scala 41:22]
  reg [21:0] mem_104; // @[RAM.scala 41:22]
  reg [21:0] mem_105; // @[RAM.scala 41:22]
  reg [21:0] mem_106; // @[RAM.scala 41:22]
  reg [21:0] mem_107; // @[RAM.scala 41:22]
  reg [21:0] mem_108; // @[RAM.scala 41:22]
  reg [21:0] mem_109; // @[RAM.scala 41:22]
  reg [21:0] mem_110; // @[RAM.scala 41:22]
  reg [21:0] mem_111; // @[RAM.scala 41:22]
  reg [21:0] mem_112; // @[RAM.scala 41:22]
  reg [21:0] mem_113; // @[RAM.scala 41:22]
  reg [21:0] mem_114; // @[RAM.scala 41:22]
  reg [21:0] mem_115; // @[RAM.scala 41:22]
  reg [21:0] mem_116; // @[RAM.scala 41:22]
  reg [21:0] mem_117; // @[RAM.scala 41:22]
  reg [21:0] mem_118; // @[RAM.scala 41:22]
  reg [21:0] mem_119; // @[RAM.scala 41:22]
  reg [21:0] mem_120; // @[RAM.scala 41:22]
  reg [21:0] mem_121; // @[RAM.scala 41:22]
  reg [21:0] mem_122; // @[RAM.scala 41:22]
  reg [21:0] mem_123; // @[RAM.scala 41:22]
  reg [21:0] mem_124; // @[RAM.scala 41:22]
  reg [21:0] mem_125; // @[RAM.scala 41:22]
  reg [21:0] mem_126; // @[RAM.scala 41:22]
  reg [21:0] mem_127; // @[RAM.scala 41:22]
  reg [21:0] mem_128; // @[RAM.scala 41:22]
  reg [21:0] mem_129; // @[RAM.scala 41:22]
  reg [21:0] mem_130; // @[RAM.scala 41:22]
  reg [21:0] mem_131; // @[RAM.scala 41:22]
  reg [21:0] mem_132; // @[RAM.scala 41:22]
  reg [21:0] mem_133; // @[RAM.scala 41:22]
  reg [21:0] mem_134; // @[RAM.scala 41:22]
  reg [21:0] mem_135; // @[RAM.scala 41:22]
  reg [21:0] mem_136; // @[RAM.scala 41:22]
  reg [21:0] mem_137; // @[RAM.scala 41:22]
  reg [21:0] mem_138; // @[RAM.scala 41:22]
  reg [21:0] mem_139; // @[RAM.scala 41:22]
  reg [21:0] mem_140; // @[RAM.scala 41:22]
  reg [21:0] mem_141; // @[RAM.scala 41:22]
  reg [21:0] mem_142; // @[RAM.scala 41:22]
  reg [21:0] mem_143; // @[RAM.scala 41:22]
  reg [21:0] mem_144; // @[RAM.scala 41:22]
  reg [21:0] mem_145; // @[RAM.scala 41:22]
  reg [21:0] mem_146; // @[RAM.scala 41:22]
  reg [21:0] mem_147; // @[RAM.scala 41:22]
  reg [21:0] mem_148; // @[RAM.scala 41:22]
  reg [21:0] mem_149; // @[RAM.scala 41:22]
  reg [21:0] mem_150; // @[RAM.scala 41:22]
  reg [21:0] mem_151; // @[RAM.scala 41:22]
  reg [21:0] mem_152; // @[RAM.scala 41:22]
  reg [21:0] mem_153; // @[RAM.scala 41:22]
  reg [21:0] mem_154; // @[RAM.scala 41:22]
  reg [21:0] mem_155; // @[RAM.scala 41:22]
  reg [21:0] mem_156; // @[RAM.scala 41:22]
  reg [21:0] mem_157; // @[RAM.scala 41:22]
  reg [21:0] mem_158; // @[RAM.scala 41:22]
  reg [21:0] mem_159; // @[RAM.scala 41:22]
  reg [21:0] mem_160; // @[RAM.scala 41:22]
  reg [21:0] mem_161; // @[RAM.scala 41:22]
  reg [21:0] mem_162; // @[RAM.scala 41:22]
  reg [21:0] mem_163; // @[RAM.scala 41:22]
  reg [21:0] mem_164; // @[RAM.scala 41:22]
  reg [21:0] mem_165; // @[RAM.scala 41:22]
  reg [21:0] mem_166; // @[RAM.scala 41:22]
  reg [21:0] mem_167; // @[RAM.scala 41:22]
  reg [21:0] mem_168; // @[RAM.scala 41:22]
  reg [21:0] mem_169; // @[RAM.scala 41:22]
  reg [21:0] mem_170; // @[RAM.scala 41:22]
  reg [21:0] mem_171; // @[RAM.scala 41:22]
  reg [21:0] mem_172; // @[RAM.scala 41:22]
  reg [21:0] mem_173; // @[RAM.scala 41:22]
  reg [21:0] mem_174; // @[RAM.scala 41:22]
  reg [21:0] mem_175; // @[RAM.scala 41:22]
  reg [21:0] mem_176; // @[RAM.scala 41:22]
  reg [21:0] mem_177; // @[RAM.scala 41:22]
  reg [21:0] mem_178; // @[RAM.scala 41:22]
  reg [21:0] mem_179; // @[RAM.scala 41:22]
  reg [21:0] mem_180; // @[RAM.scala 41:22]
  reg [21:0] mem_181; // @[RAM.scala 41:22]
  reg [21:0] mem_182; // @[RAM.scala 41:22]
  reg [21:0] mem_183; // @[RAM.scala 41:22]
  reg [21:0] mem_184; // @[RAM.scala 41:22]
  reg [21:0] mem_185; // @[RAM.scala 41:22]
  reg [21:0] mem_186; // @[RAM.scala 41:22]
  reg [21:0] mem_187; // @[RAM.scala 41:22]
  reg [21:0] mem_188; // @[RAM.scala 41:22]
  reg [21:0] mem_189; // @[RAM.scala 41:22]
  reg [21:0] mem_190; // @[RAM.scala 41:22]
  reg [21:0] mem_191; // @[RAM.scala 41:22]
  reg [21:0] mem_192; // @[RAM.scala 41:22]
  reg [21:0] mem_193; // @[RAM.scala 41:22]
  reg [21:0] mem_194; // @[RAM.scala 41:22]
  reg [21:0] mem_195; // @[RAM.scala 41:22]
  reg [21:0] mem_196; // @[RAM.scala 41:22]
  reg [21:0] mem_197; // @[RAM.scala 41:22]
  reg [21:0] mem_198; // @[RAM.scala 41:22]
  reg [21:0] mem_199; // @[RAM.scala 41:22]
  reg [21:0] mem_200; // @[RAM.scala 41:22]
  reg [21:0] mem_201; // @[RAM.scala 41:22]
  reg [21:0] mem_202; // @[RAM.scala 41:22]
  reg [21:0] mem_203; // @[RAM.scala 41:22]
  reg [21:0] mem_204; // @[RAM.scala 41:22]
  reg [21:0] mem_205; // @[RAM.scala 41:22]
  reg [21:0] mem_206; // @[RAM.scala 41:22]
  reg [21:0] mem_207; // @[RAM.scala 41:22]
  reg [21:0] mem_208; // @[RAM.scala 41:22]
  reg [21:0] mem_209; // @[RAM.scala 41:22]
  reg [21:0] mem_210; // @[RAM.scala 41:22]
  reg [21:0] mem_211; // @[RAM.scala 41:22]
  reg [21:0] mem_212; // @[RAM.scala 41:22]
  reg [21:0] mem_213; // @[RAM.scala 41:22]
  reg [21:0] mem_214; // @[RAM.scala 41:22]
  reg [21:0] mem_215; // @[RAM.scala 41:22]
  reg [21:0] mem_216; // @[RAM.scala 41:22]
  reg [21:0] mem_217; // @[RAM.scala 41:22]
  reg [21:0] mem_218; // @[RAM.scala 41:22]
  reg [21:0] mem_219; // @[RAM.scala 41:22]
  reg [21:0] mem_220; // @[RAM.scala 41:22]
  reg [21:0] mem_221; // @[RAM.scala 41:22]
  reg [21:0] mem_222; // @[RAM.scala 41:22]
  reg [21:0] mem_223; // @[RAM.scala 41:22]
  reg [21:0] mem_224; // @[RAM.scala 41:22]
  reg [21:0] mem_225; // @[RAM.scala 41:22]
  reg [21:0] mem_226; // @[RAM.scala 41:22]
  reg [21:0] mem_227; // @[RAM.scala 41:22]
  reg [21:0] mem_228; // @[RAM.scala 41:22]
  reg [21:0] mem_229; // @[RAM.scala 41:22]
  reg [21:0] mem_230; // @[RAM.scala 41:22]
  reg [21:0] mem_231; // @[RAM.scala 41:22]
  reg [21:0] mem_232; // @[RAM.scala 41:22]
  reg [21:0] mem_233; // @[RAM.scala 41:22]
  reg [21:0] mem_234; // @[RAM.scala 41:22]
  reg [21:0] mem_235; // @[RAM.scala 41:22]
  reg [21:0] mem_236; // @[RAM.scala 41:22]
  reg [21:0] mem_237; // @[RAM.scala 41:22]
  reg [21:0] mem_238; // @[RAM.scala 41:22]
  reg [21:0] mem_239; // @[RAM.scala 41:22]
  reg [21:0] mem_240; // @[RAM.scala 41:22]
  reg [21:0] mem_241; // @[RAM.scala 41:22]
  reg [21:0] mem_242; // @[RAM.scala 41:22]
  reg [21:0] mem_243; // @[RAM.scala 41:22]
  reg [21:0] mem_244; // @[RAM.scala 41:22]
  reg [21:0] mem_245; // @[RAM.scala 41:22]
  reg [21:0] mem_246; // @[RAM.scala 41:22]
  reg [21:0] mem_247; // @[RAM.scala 41:22]
  reg [21:0] mem_248; // @[RAM.scala 41:22]
  reg [21:0] mem_249; // @[RAM.scala 41:22]
  reg [21:0] mem_250; // @[RAM.scala 41:22]
  reg [21:0] mem_251; // @[RAM.scala 41:22]
  reg [21:0] mem_252; // @[RAM.scala 41:22]
  reg [21:0] mem_253; // @[RAM.scala 41:22]
  reg [21:0] mem_254; // @[RAM.scala 41:22]
  reg [21:0] mem_255; // @[RAM.scala 41:22]
  reg [21:0] io_douta_REG; // @[RAM.scala 43:24]
  wire [21:0] _GEN_1 = 8'h1 == io_addra ? mem_1 : mem_0; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_2 = 8'h2 == io_addra ? mem_2 : _GEN_1; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_3 = 8'h3 == io_addra ? mem_3 : _GEN_2; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_4 = 8'h4 == io_addra ? mem_4 : _GEN_3; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_5 = 8'h5 == io_addra ? mem_5 : _GEN_4; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_6 = 8'h6 == io_addra ? mem_6 : _GEN_5; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_7 = 8'h7 == io_addra ? mem_7 : _GEN_6; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_8 = 8'h8 == io_addra ? mem_8 : _GEN_7; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_9 = 8'h9 == io_addra ? mem_9 : _GEN_8; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_10 = 8'ha == io_addra ? mem_10 : _GEN_9; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_11 = 8'hb == io_addra ? mem_11 : _GEN_10; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_12 = 8'hc == io_addra ? mem_12 : _GEN_11; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_13 = 8'hd == io_addra ? mem_13 : _GEN_12; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_14 = 8'he == io_addra ? mem_14 : _GEN_13; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_15 = 8'hf == io_addra ? mem_15 : _GEN_14; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_16 = 8'h10 == io_addra ? mem_16 : _GEN_15; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_17 = 8'h11 == io_addra ? mem_17 : _GEN_16; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_18 = 8'h12 == io_addra ? mem_18 : _GEN_17; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_19 = 8'h13 == io_addra ? mem_19 : _GEN_18; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_20 = 8'h14 == io_addra ? mem_20 : _GEN_19; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_21 = 8'h15 == io_addra ? mem_21 : _GEN_20; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_22 = 8'h16 == io_addra ? mem_22 : _GEN_21; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_23 = 8'h17 == io_addra ? mem_23 : _GEN_22; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_24 = 8'h18 == io_addra ? mem_24 : _GEN_23; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_25 = 8'h19 == io_addra ? mem_25 : _GEN_24; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_26 = 8'h1a == io_addra ? mem_26 : _GEN_25; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_27 = 8'h1b == io_addra ? mem_27 : _GEN_26; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_28 = 8'h1c == io_addra ? mem_28 : _GEN_27; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_29 = 8'h1d == io_addra ? mem_29 : _GEN_28; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_30 = 8'h1e == io_addra ? mem_30 : _GEN_29; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_31 = 8'h1f == io_addra ? mem_31 : _GEN_30; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_32 = 8'h20 == io_addra ? mem_32 : _GEN_31; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_33 = 8'h21 == io_addra ? mem_33 : _GEN_32; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_34 = 8'h22 == io_addra ? mem_34 : _GEN_33; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_35 = 8'h23 == io_addra ? mem_35 : _GEN_34; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_36 = 8'h24 == io_addra ? mem_36 : _GEN_35; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_37 = 8'h25 == io_addra ? mem_37 : _GEN_36; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_38 = 8'h26 == io_addra ? mem_38 : _GEN_37; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_39 = 8'h27 == io_addra ? mem_39 : _GEN_38; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_40 = 8'h28 == io_addra ? mem_40 : _GEN_39; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_41 = 8'h29 == io_addra ? mem_41 : _GEN_40; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_42 = 8'h2a == io_addra ? mem_42 : _GEN_41; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_43 = 8'h2b == io_addra ? mem_43 : _GEN_42; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_44 = 8'h2c == io_addra ? mem_44 : _GEN_43; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_45 = 8'h2d == io_addra ? mem_45 : _GEN_44; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_46 = 8'h2e == io_addra ? mem_46 : _GEN_45; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_47 = 8'h2f == io_addra ? mem_47 : _GEN_46; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_48 = 8'h30 == io_addra ? mem_48 : _GEN_47; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_49 = 8'h31 == io_addra ? mem_49 : _GEN_48; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_50 = 8'h32 == io_addra ? mem_50 : _GEN_49; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_51 = 8'h33 == io_addra ? mem_51 : _GEN_50; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_52 = 8'h34 == io_addra ? mem_52 : _GEN_51; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_53 = 8'h35 == io_addra ? mem_53 : _GEN_52; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_54 = 8'h36 == io_addra ? mem_54 : _GEN_53; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_55 = 8'h37 == io_addra ? mem_55 : _GEN_54; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_56 = 8'h38 == io_addra ? mem_56 : _GEN_55; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_57 = 8'h39 == io_addra ? mem_57 : _GEN_56; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_58 = 8'h3a == io_addra ? mem_58 : _GEN_57; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_59 = 8'h3b == io_addra ? mem_59 : _GEN_58; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_60 = 8'h3c == io_addra ? mem_60 : _GEN_59; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_61 = 8'h3d == io_addra ? mem_61 : _GEN_60; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_62 = 8'h3e == io_addra ? mem_62 : _GEN_61; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_63 = 8'h3f == io_addra ? mem_63 : _GEN_62; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_64 = 8'h40 == io_addra ? mem_64 : _GEN_63; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_65 = 8'h41 == io_addra ? mem_65 : _GEN_64; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_66 = 8'h42 == io_addra ? mem_66 : _GEN_65; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_67 = 8'h43 == io_addra ? mem_67 : _GEN_66; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_68 = 8'h44 == io_addra ? mem_68 : _GEN_67; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_69 = 8'h45 == io_addra ? mem_69 : _GEN_68; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_70 = 8'h46 == io_addra ? mem_70 : _GEN_69; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_71 = 8'h47 == io_addra ? mem_71 : _GEN_70; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_72 = 8'h48 == io_addra ? mem_72 : _GEN_71; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_73 = 8'h49 == io_addra ? mem_73 : _GEN_72; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_74 = 8'h4a == io_addra ? mem_74 : _GEN_73; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_75 = 8'h4b == io_addra ? mem_75 : _GEN_74; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_76 = 8'h4c == io_addra ? mem_76 : _GEN_75; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_77 = 8'h4d == io_addra ? mem_77 : _GEN_76; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_78 = 8'h4e == io_addra ? mem_78 : _GEN_77; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_79 = 8'h4f == io_addra ? mem_79 : _GEN_78; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_80 = 8'h50 == io_addra ? mem_80 : _GEN_79; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_81 = 8'h51 == io_addra ? mem_81 : _GEN_80; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_82 = 8'h52 == io_addra ? mem_82 : _GEN_81; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_83 = 8'h53 == io_addra ? mem_83 : _GEN_82; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_84 = 8'h54 == io_addra ? mem_84 : _GEN_83; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_85 = 8'h55 == io_addra ? mem_85 : _GEN_84; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_86 = 8'h56 == io_addra ? mem_86 : _GEN_85; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_87 = 8'h57 == io_addra ? mem_87 : _GEN_86; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_88 = 8'h58 == io_addra ? mem_88 : _GEN_87; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_89 = 8'h59 == io_addra ? mem_89 : _GEN_88; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_90 = 8'h5a == io_addra ? mem_90 : _GEN_89; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_91 = 8'h5b == io_addra ? mem_91 : _GEN_90; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_92 = 8'h5c == io_addra ? mem_92 : _GEN_91; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_93 = 8'h5d == io_addra ? mem_93 : _GEN_92; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_94 = 8'h5e == io_addra ? mem_94 : _GEN_93; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_95 = 8'h5f == io_addra ? mem_95 : _GEN_94; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_96 = 8'h60 == io_addra ? mem_96 : _GEN_95; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_97 = 8'h61 == io_addra ? mem_97 : _GEN_96; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_98 = 8'h62 == io_addra ? mem_98 : _GEN_97; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_99 = 8'h63 == io_addra ? mem_99 : _GEN_98; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_100 = 8'h64 == io_addra ? mem_100 : _GEN_99; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_101 = 8'h65 == io_addra ? mem_101 : _GEN_100; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_102 = 8'h66 == io_addra ? mem_102 : _GEN_101; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_103 = 8'h67 == io_addra ? mem_103 : _GEN_102; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_104 = 8'h68 == io_addra ? mem_104 : _GEN_103; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_105 = 8'h69 == io_addra ? mem_105 : _GEN_104; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_106 = 8'h6a == io_addra ? mem_106 : _GEN_105; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_107 = 8'h6b == io_addra ? mem_107 : _GEN_106; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_108 = 8'h6c == io_addra ? mem_108 : _GEN_107; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_109 = 8'h6d == io_addra ? mem_109 : _GEN_108; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_110 = 8'h6e == io_addra ? mem_110 : _GEN_109; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_111 = 8'h6f == io_addra ? mem_111 : _GEN_110; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_112 = 8'h70 == io_addra ? mem_112 : _GEN_111; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_113 = 8'h71 == io_addra ? mem_113 : _GEN_112; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_114 = 8'h72 == io_addra ? mem_114 : _GEN_113; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_115 = 8'h73 == io_addra ? mem_115 : _GEN_114; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_116 = 8'h74 == io_addra ? mem_116 : _GEN_115; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_117 = 8'h75 == io_addra ? mem_117 : _GEN_116; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_118 = 8'h76 == io_addra ? mem_118 : _GEN_117; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_119 = 8'h77 == io_addra ? mem_119 : _GEN_118; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_120 = 8'h78 == io_addra ? mem_120 : _GEN_119; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_121 = 8'h79 == io_addra ? mem_121 : _GEN_120; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_122 = 8'h7a == io_addra ? mem_122 : _GEN_121; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_123 = 8'h7b == io_addra ? mem_123 : _GEN_122; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_124 = 8'h7c == io_addra ? mem_124 : _GEN_123; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_125 = 8'h7d == io_addra ? mem_125 : _GEN_124; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_126 = 8'h7e == io_addra ? mem_126 : _GEN_125; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_127 = 8'h7f == io_addra ? mem_127 : _GEN_126; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_128 = 8'h80 == io_addra ? mem_128 : _GEN_127; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_129 = 8'h81 == io_addra ? mem_129 : _GEN_128; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_130 = 8'h82 == io_addra ? mem_130 : _GEN_129; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_131 = 8'h83 == io_addra ? mem_131 : _GEN_130; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_132 = 8'h84 == io_addra ? mem_132 : _GEN_131; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_133 = 8'h85 == io_addra ? mem_133 : _GEN_132; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_134 = 8'h86 == io_addra ? mem_134 : _GEN_133; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_135 = 8'h87 == io_addra ? mem_135 : _GEN_134; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_136 = 8'h88 == io_addra ? mem_136 : _GEN_135; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_137 = 8'h89 == io_addra ? mem_137 : _GEN_136; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_138 = 8'h8a == io_addra ? mem_138 : _GEN_137; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_139 = 8'h8b == io_addra ? mem_139 : _GEN_138; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_140 = 8'h8c == io_addra ? mem_140 : _GEN_139; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_141 = 8'h8d == io_addra ? mem_141 : _GEN_140; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_142 = 8'h8e == io_addra ? mem_142 : _GEN_141; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_143 = 8'h8f == io_addra ? mem_143 : _GEN_142; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_144 = 8'h90 == io_addra ? mem_144 : _GEN_143; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_145 = 8'h91 == io_addra ? mem_145 : _GEN_144; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_146 = 8'h92 == io_addra ? mem_146 : _GEN_145; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_147 = 8'h93 == io_addra ? mem_147 : _GEN_146; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_148 = 8'h94 == io_addra ? mem_148 : _GEN_147; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_149 = 8'h95 == io_addra ? mem_149 : _GEN_148; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_150 = 8'h96 == io_addra ? mem_150 : _GEN_149; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_151 = 8'h97 == io_addra ? mem_151 : _GEN_150; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_152 = 8'h98 == io_addra ? mem_152 : _GEN_151; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_153 = 8'h99 == io_addra ? mem_153 : _GEN_152; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_154 = 8'h9a == io_addra ? mem_154 : _GEN_153; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_155 = 8'h9b == io_addra ? mem_155 : _GEN_154; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_156 = 8'h9c == io_addra ? mem_156 : _GEN_155; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_157 = 8'h9d == io_addra ? mem_157 : _GEN_156; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_158 = 8'h9e == io_addra ? mem_158 : _GEN_157; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_159 = 8'h9f == io_addra ? mem_159 : _GEN_158; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_160 = 8'ha0 == io_addra ? mem_160 : _GEN_159; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_161 = 8'ha1 == io_addra ? mem_161 : _GEN_160; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_162 = 8'ha2 == io_addra ? mem_162 : _GEN_161; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_163 = 8'ha3 == io_addra ? mem_163 : _GEN_162; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_164 = 8'ha4 == io_addra ? mem_164 : _GEN_163; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_165 = 8'ha5 == io_addra ? mem_165 : _GEN_164; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_166 = 8'ha6 == io_addra ? mem_166 : _GEN_165; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_167 = 8'ha7 == io_addra ? mem_167 : _GEN_166; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_168 = 8'ha8 == io_addra ? mem_168 : _GEN_167; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_169 = 8'ha9 == io_addra ? mem_169 : _GEN_168; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_170 = 8'haa == io_addra ? mem_170 : _GEN_169; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_171 = 8'hab == io_addra ? mem_171 : _GEN_170; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_172 = 8'hac == io_addra ? mem_172 : _GEN_171; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_173 = 8'had == io_addra ? mem_173 : _GEN_172; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_174 = 8'hae == io_addra ? mem_174 : _GEN_173; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_175 = 8'haf == io_addra ? mem_175 : _GEN_174; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_176 = 8'hb0 == io_addra ? mem_176 : _GEN_175; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_177 = 8'hb1 == io_addra ? mem_177 : _GEN_176; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_178 = 8'hb2 == io_addra ? mem_178 : _GEN_177; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_179 = 8'hb3 == io_addra ? mem_179 : _GEN_178; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_180 = 8'hb4 == io_addra ? mem_180 : _GEN_179; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_181 = 8'hb5 == io_addra ? mem_181 : _GEN_180; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_182 = 8'hb6 == io_addra ? mem_182 : _GEN_181; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_183 = 8'hb7 == io_addra ? mem_183 : _GEN_182; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_184 = 8'hb8 == io_addra ? mem_184 : _GEN_183; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_185 = 8'hb9 == io_addra ? mem_185 : _GEN_184; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_186 = 8'hba == io_addra ? mem_186 : _GEN_185; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_187 = 8'hbb == io_addra ? mem_187 : _GEN_186; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_188 = 8'hbc == io_addra ? mem_188 : _GEN_187; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_189 = 8'hbd == io_addra ? mem_189 : _GEN_188; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_190 = 8'hbe == io_addra ? mem_190 : _GEN_189; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_191 = 8'hbf == io_addra ? mem_191 : _GEN_190; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_192 = 8'hc0 == io_addra ? mem_192 : _GEN_191; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_193 = 8'hc1 == io_addra ? mem_193 : _GEN_192; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_194 = 8'hc2 == io_addra ? mem_194 : _GEN_193; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_195 = 8'hc3 == io_addra ? mem_195 : _GEN_194; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_196 = 8'hc4 == io_addra ? mem_196 : _GEN_195; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_197 = 8'hc5 == io_addra ? mem_197 : _GEN_196; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_198 = 8'hc6 == io_addra ? mem_198 : _GEN_197; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_199 = 8'hc7 == io_addra ? mem_199 : _GEN_198; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_200 = 8'hc8 == io_addra ? mem_200 : _GEN_199; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_201 = 8'hc9 == io_addra ? mem_201 : _GEN_200; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_202 = 8'hca == io_addra ? mem_202 : _GEN_201; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_203 = 8'hcb == io_addra ? mem_203 : _GEN_202; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_204 = 8'hcc == io_addra ? mem_204 : _GEN_203; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_205 = 8'hcd == io_addra ? mem_205 : _GEN_204; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_206 = 8'hce == io_addra ? mem_206 : _GEN_205; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_207 = 8'hcf == io_addra ? mem_207 : _GEN_206; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_208 = 8'hd0 == io_addra ? mem_208 : _GEN_207; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_209 = 8'hd1 == io_addra ? mem_209 : _GEN_208; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_210 = 8'hd2 == io_addra ? mem_210 : _GEN_209; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_211 = 8'hd3 == io_addra ? mem_211 : _GEN_210; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_212 = 8'hd4 == io_addra ? mem_212 : _GEN_211; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_213 = 8'hd5 == io_addra ? mem_213 : _GEN_212; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_214 = 8'hd6 == io_addra ? mem_214 : _GEN_213; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_215 = 8'hd7 == io_addra ? mem_215 : _GEN_214; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_216 = 8'hd8 == io_addra ? mem_216 : _GEN_215; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_217 = 8'hd9 == io_addra ? mem_217 : _GEN_216; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_218 = 8'hda == io_addra ? mem_218 : _GEN_217; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_219 = 8'hdb == io_addra ? mem_219 : _GEN_218; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_220 = 8'hdc == io_addra ? mem_220 : _GEN_219; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_221 = 8'hdd == io_addra ? mem_221 : _GEN_220; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_222 = 8'hde == io_addra ? mem_222 : _GEN_221; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_223 = 8'hdf == io_addra ? mem_223 : _GEN_222; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_224 = 8'he0 == io_addra ? mem_224 : _GEN_223; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_225 = 8'he1 == io_addra ? mem_225 : _GEN_224; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_226 = 8'he2 == io_addra ? mem_226 : _GEN_225; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_227 = 8'he3 == io_addra ? mem_227 : _GEN_226; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_228 = 8'he4 == io_addra ? mem_228 : _GEN_227; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_229 = 8'he5 == io_addra ? mem_229 : _GEN_228; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_230 = 8'he6 == io_addra ? mem_230 : _GEN_229; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_231 = 8'he7 == io_addra ? mem_231 : _GEN_230; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_232 = 8'he8 == io_addra ? mem_232 : _GEN_231; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_233 = 8'he9 == io_addra ? mem_233 : _GEN_232; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_234 = 8'hea == io_addra ? mem_234 : _GEN_233; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_235 = 8'heb == io_addra ? mem_235 : _GEN_234; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_236 = 8'hec == io_addra ? mem_236 : _GEN_235; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_237 = 8'hed == io_addra ? mem_237 : _GEN_236; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_238 = 8'hee == io_addra ? mem_238 : _GEN_237; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_239 = 8'hef == io_addra ? mem_239 : _GEN_238; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_240 = 8'hf0 == io_addra ? mem_240 : _GEN_239; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_241 = 8'hf1 == io_addra ? mem_241 : _GEN_240; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_242 = 8'hf2 == io_addra ? mem_242 : _GEN_241; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_243 = 8'hf3 == io_addra ? mem_243 : _GEN_242; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_244 = 8'hf4 == io_addra ? mem_244 : _GEN_243; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_245 = 8'hf5 == io_addra ? mem_245 : _GEN_244; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_246 = 8'hf6 == io_addra ? mem_246 : _GEN_245; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_247 = 8'hf7 == io_addra ? mem_247 : _GEN_246; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_248 = 8'hf8 == io_addra ? mem_248 : _GEN_247; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_249 = 8'hf9 == io_addra ? mem_249 : _GEN_248; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_250 = 8'hfa == io_addra ? mem_250 : _GEN_249; // @[RAM.scala 43:24 RAM.scala 43:24]
  wire [21:0] _GEN_251 = 8'hfb == io_addra ? mem_251 : _GEN_250; // @[RAM.scala 43:24 RAM.scala 43:24]
  assign io_douta = io_douta_REG; // @[RAM.scala 43:14]
  always @(posedge clock) begin
    if (reset) begin // @[RAM.scala 41:22]
      mem_0 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h0 == io_addrb) begin // @[RAM.scala 50:23]
        mem_0 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_1 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h1 == io_addrb) begin // @[RAM.scala 50:23]
        mem_1 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_2 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h2 == io_addrb) begin // @[RAM.scala 50:23]
        mem_2 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_3 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h3 == io_addrb) begin // @[RAM.scala 50:23]
        mem_3 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_4 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h4 == io_addrb) begin // @[RAM.scala 50:23]
        mem_4 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_5 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h5 == io_addrb) begin // @[RAM.scala 50:23]
        mem_5 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_6 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h6 == io_addrb) begin // @[RAM.scala 50:23]
        mem_6 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_7 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h7 == io_addrb) begin // @[RAM.scala 50:23]
        mem_7 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_8 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h8 == io_addrb) begin // @[RAM.scala 50:23]
        mem_8 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_9 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h9 == io_addrb) begin // @[RAM.scala 50:23]
        mem_9 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_10 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha == io_addrb) begin // @[RAM.scala 50:23]
        mem_10 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_11 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb == io_addrb) begin // @[RAM.scala 50:23]
        mem_11 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_12 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc == io_addrb) begin // @[RAM.scala 50:23]
        mem_12 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_13 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd == io_addrb) begin // @[RAM.scala 50:23]
        mem_13 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_14 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he == io_addrb) begin // @[RAM.scala 50:23]
        mem_14 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_15 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf == io_addrb) begin // @[RAM.scala 50:23]
        mem_15 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_16 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h10 == io_addrb) begin // @[RAM.scala 50:23]
        mem_16 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_17 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h11 == io_addrb) begin // @[RAM.scala 50:23]
        mem_17 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_18 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h12 == io_addrb) begin // @[RAM.scala 50:23]
        mem_18 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_19 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h13 == io_addrb) begin // @[RAM.scala 50:23]
        mem_19 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_20 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h14 == io_addrb) begin // @[RAM.scala 50:23]
        mem_20 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_21 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h15 == io_addrb) begin // @[RAM.scala 50:23]
        mem_21 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_22 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h16 == io_addrb) begin // @[RAM.scala 50:23]
        mem_22 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_23 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h17 == io_addrb) begin // @[RAM.scala 50:23]
        mem_23 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_24 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h18 == io_addrb) begin // @[RAM.scala 50:23]
        mem_24 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_25 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h19 == io_addrb) begin // @[RAM.scala 50:23]
        mem_25 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_26 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h1a == io_addrb) begin // @[RAM.scala 50:23]
        mem_26 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_27 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h1b == io_addrb) begin // @[RAM.scala 50:23]
        mem_27 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_28 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h1c == io_addrb) begin // @[RAM.scala 50:23]
        mem_28 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_29 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h1d == io_addrb) begin // @[RAM.scala 50:23]
        mem_29 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_30 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h1e == io_addrb) begin // @[RAM.scala 50:23]
        mem_30 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_31 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h1f == io_addrb) begin // @[RAM.scala 50:23]
        mem_31 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_32 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h20 == io_addrb) begin // @[RAM.scala 50:23]
        mem_32 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_33 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h21 == io_addrb) begin // @[RAM.scala 50:23]
        mem_33 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_34 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h22 == io_addrb) begin // @[RAM.scala 50:23]
        mem_34 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_35 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h23 == io_addrb) begin // @[RAM.scala 50:23]
        mem_35 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_36 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h24 == io_addrb) begin // @[RAM.scala 50:23]
        mem_36 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_37 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h25 == io_addrb) begin // @[RAM.scala 50:23]
        mem_37 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_38 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h26 == io_addrb) begin // @[RAM.scala 50:23]
        mem_38 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_39 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h27 == io_addrb) begin // @[RAM.scala 50:23]
        mem_39 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_40 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h28 == io_addrb) begin // @[RAM.scala 50:23]
        mem_40 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_41 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h29 == io_addrb) begin // @[RAM.scala 50:23]
        mem_41 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_42 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h2a == io_addrb) begin // @[RAM.scala 50:23]
        mem_42 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_43 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h2b == io_addrb) begin // @[RAM.scala 50:23]
        mem_43 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_44 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h2c == io_addrb) begin // @[RAM.scala 50:23]
        mem_44 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_45 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h2d == io_addrb) begin // @[RAM.scala 50:23]
        mem_45 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_46 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h2e == io_addrb) begin // @[RAM.scala 50:23]
        mem_46 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_47 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h2f == io_addrb) begin // @[RAM.scala 50:23]
        mem_47 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_48 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h30 == io_addrb) begin // @[RAM.scala 50:23]
        mem_48 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_49 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h31 == io_addrb) begin // @[RAM.scala 50:23]
        mem_49 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_50 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h32 == io_addrb) begin // @[RAM.scala 50:23]
        mem_50 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_51 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h33 == io_addrb) begin // @[RAM.scala 50:23]
        mem_51 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_52 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h34 == io_addrb) begin // @[RAM.scala 50:23]
        mem_52 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_53 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h35 == io_addrb) begin // @[RAM.scala 50:23]
        mem_53 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_54 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h36 == io_addrb) begin // @[RAM.scala 50:23]
        mem_54 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_55 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h37 == io_addrb) begin // @[RAM.scala 50:23]
        mem_55 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_56 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h38 == io_addrb) begin // @[RAM.scala 50:23]
        mem_56 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_57 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h39 == io_addrb) begin // @[RAM.scala 50:23]
        mem_57 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_58 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h3a == io_addrb) begin // @[RAM.scala 50:23]
        mem_58 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_59 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h3b == io_addrb) begin // @[RAM.scala 50:23]
        mem_59 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_60 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h3c == io_addrb) begin // @[RAM.scala 50:23]
        mem_60 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_61 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h3d == io_addrb) begin // @[RAM.scala 50:23]
        mem_61 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_62 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h3e == io_addrb) begin // @[RAM.scala 50:23]
        mem_62 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_63 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h3f == io_addrb) begin // @[RAM.scala 50:23]
        mem_63 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_64 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h40 == io_addrb) begin // @[RAM.scala 50:23]
        mem_64 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_65 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h41 == io_addrb) begin // @[RAM.scala 50:23]
        mem_65 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_66 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h42 == io_addrb) begin // @[RAM.scala 50:23]
        mem_66 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_67 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h43 == io_addrb) begin // @[RAM.scala 50:23]
        mem_67 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_68 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h44 == io_addrb) begin // @[RAM.scala 50:23]
        mem_68 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_69 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h45 == io_addrb) begin // @[RAM.scala 50:23]
        mem_69 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_70 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h46 == io_addrb) begin // @[RAM.scala 50:23]
        mem_70 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_71 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h47 == io_addrb) begin // @[RAM.scala 50:23]
        mem_71 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_72 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h48 == io_addrb) begin // @[RAM.scala 50:23]
        mem_72 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_73 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h49 == io_addrb) begin // @[RAM.scala 50:23]
        mem_73 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_74 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h4a == io_addrb) begin // @[RAM.scala 50:23]
        mem_74 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_75 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h4b == io_addrb) begin // @[RAM.scala 50:23]
        mem_75 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_76 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h4c == io_addrb) begin // @[RAM.scala 50:23]
        mem_76 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_77 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h4d == io_addrb) begin // @[RAM.scala 50:23]
        mem_77 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_78 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h4e == io_addrb) begin // @[RAM.scala 50:23]
        mem_78 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_79 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h4f == io_addrb) begin // @[RAM.scala 50:23]
        mem_79 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_80 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h50 == io_addrb) begin // @[RAM.scala 50:23]
        mem_80 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_81 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h51 == io_addrb) begin // @[RAM.scala 50:23]
        mem_81 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_82 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h52 == io_addrb) begin // @[RAM.scala 50:23]
        mem_82 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_83 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h53 == io_addrb) begin // @[RAM.scala 50:23]
        mem_83 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_84 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h54 == io_addrb) begin // @[RAM.scala 50:23]
        mem_84 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_85 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h55 == io_addrb) begin // @[RAM.scala 50:23]
        mem_85 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_86 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h56 == io_addrb) begin // @[RAM.scala 50:23]
        mem_86 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_87 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h57 == io_addrb) begin // @[RAM.scala 50:23]
        mem_87 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_88 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h58 == io_addrb) begin // @[RAM.scala 50:23]
        mem_88 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_89 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h59 == io_addrb) begin // @[RAM.scala 50:23]
        mem_89 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_90 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h5a == io_addrb) begin // @[RAM.scala 50:23]
        mem_90 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_91 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h5b == io_addrb) begin // @[RAM.scala 50:23]
        mem_91 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_92 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h5c == io_addrb) begin // @[RAM.scala 50:23]
        mem_92 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_93 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h5d == io_addrb) begin // @[RAM.scala 50:23]
        mem_93 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_94 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h5e == io_addrb) begin // @[RAM.scala 50:23]
        mem_94 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_95 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h5f == io_addrb) begin // @[RAM.scala 50:23]
        mem_95 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_96 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h60 == io_addrb) begin // @[RAM.scala 50:23]
        mem_96 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_97 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h61 == io_addrb) begin // @[RAM.scala 50:23]
        mem_97 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_98 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h62 == io_addrb) begin // @[RAM.scala 50:23]
        mem_98 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_99 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h63 == io_addrb) begin // @[RAM.scala 50:23]
        mem_99 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_100 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h64 == io_addrb) begin // @[RAM.scala 50:23]
        mem_100 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_101 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h65 == io_addrb) begin // @[RAM.scala 50:23]
        mem_101 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_102 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h66 == io_addrb) begin // @[RAM.scala 50:23]
        mem_102 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_103 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h67 == io_addrb) begin // @[RAM.scala 50:23]
        mem_103 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_104 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h68 == io_addrb) begin // @[RAM.scala 50:23]
        mem_104 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_105 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h69 == io_addrb) begin // @[RAM.scala 50:23]
        mem_105 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_106 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h6a == io_addrb) begin // @[RAM.scala 50:23]
        mem_106 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_107 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h6b == io_addrb) begin // @[RAM.scala 50:23]
        mem_107 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_108 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h6c == io_addrb) begin // @[RAM.scala 50:23]
        mem_108 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_109 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h6d == io_addrb) begin // @[RAM.scala 50:23]
        mem_109 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_110 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h6e == io_addrb) begin // @[RAM.scala 50:23]
        mem_110 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_111 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h6f == io_addrb) begin // @[RAM.scala 50:23]
        mem_111 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_112 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h70 == io_addrb) begin // @[RAM.scala 50:23]
        mem_112 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_113 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h71 == io_addrb) begin // @[RAM.scala 50:23]
        mem_113 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_114 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h72 == io_addrb) begin // @[RAM.scala 50:23]
        mem_114 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_115 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h73 == io_addrb) begin // @[RAM.scala 50:23]
        mem_115 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_116 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h74 == io_addrb) begin // @[RAM.scala 50:23]
        mem_116 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_117 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h75 == io_addrb) begin // @[RAM.scala 50:23]
        mem_117 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_118 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h76 == io_addrb) begin // @[RAM.scala 50:23]
        mem_118 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_119 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h77 == io_addrb) begin // @[RAM.scala 50:23]
        mem_119 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_120 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h78 == io_addrb) begin // @[RAM.scala 50:23]
        mem_120 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_121 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h79 == io_addrb) begin // @[RAM.scala 50:23]
        mem_121 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_122 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h7a == io_addrb) begin // @[RAM.scala 50:23]
        mem_122 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_123 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h7b == io_addrb) begin // @[RAM.scala 50:23]
        mem_123 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_124 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h7c == io_addrb) begin // @[RAM.scala 50:23]
        mem_124 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_125 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h7d == io_addrb) begin // @[RAM.scala 50:23]
        mem_125 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_126 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h7e == io_addrb) begin // @[RAM.scala 50:23]
        mem_126 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_127 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h7f == io_addrb) begin // @[RAM.scala 50:23]
        mem_127 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_128 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h80 == io_addrb) begin // @[RAM.scala 50:23]
        mem_128 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_129 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h81 == io_addrb) begin // @[RAM.scala 50:23]
        mem_129 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_130 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h82 == io_addrb) begin // @[RAM.scala 50:23]
        mem_130 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_131 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h83 == io_addrb) begin // @[RAM.scala 50:23]
        mem_131 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_132 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h84 == io_addrb) begin // @[RAM.scala 50:23]
        mem_132 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_133 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h85 == io_addrb) begin // @[RAM.scala 50:23]
        mem_133 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_134 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h86 == io_addrb) begin // @[RAM.scala 50:23]
        mem_134 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_135 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h87 == io_addrb) begin // @[RAM.scala 50:23]
        mem_135 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_136 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h88 == io_addrb) begin // @[RAM.scala 50:23]
        mem_136 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_137 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h89 == io_addrb) begin // @[RAM.scala 50:23]
        mem_137 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_138 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h8a == io_addrb) begin // @[RAM.scala 50:23]
        mem_138 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_139 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h8b == io_addrb) begin // @[RAM.scala 50:23]
        mem_139 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_140 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h8c == io_addrb) begin // @[RAM.scala 50:23]
        mem_140 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_141 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h8d == io_addrb) begin // @[RAM.scala 50:23]
        mem_141 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_142 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h8e == io_addrb) begin // @[RAM.scala 50:23]
        mem_142 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_143 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h8f == io_addrb) begin // @[RAM.scala 50:23]
        mem_143 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_144 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h90 == io_addrb) begin // @[RAM.scala 50:23]
        mem_144 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_145 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h91 == io_addrb) begin // @[RAM.scala 50:23]
        mem_145 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_146 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h92 == io_addrb) begin // @[RAM.scala 50:23]
        mem_146 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_147 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h93 == io_addrb) begin // @[RAM.scala 50:23]
        mem_147 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_148 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h94 == io_addrb) begin // @[RAM.scala 50:23]
        mem_148 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_149 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h95 == io_addrb) begin // @[RAM.scala 50:23]
        mem_149 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_150 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h96 == io_addrb) begin // @[RAM.scala 50:23]
        mem_150 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_151 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h97 == io_addrb) begin // @[RAM.scala 50:23]
        mem_151 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_152 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h98 == io_addrb) begin // @[RAM.scala 50:23]
        mem_152 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_153 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h99 == io_addrb) begin // @[RAM.scala 50:23]
        mem_153 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_154 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h9a == io_addrb) begin // @[RAM.scala 50:23]
        mem_154 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_155 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h9b == io_addrb) begin // @[RAM.scala 50:23]
        mem_155 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_156 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h9c == io_addrb) begin // @[RAM.scala 50:23]
        mem_156 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_157 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h9d == io_addrb) begin // @[RAM.scala 50:23]
        mem_157 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_158 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h9e == io_addrb) begin // @[RAM.scala 50:23]
        mem_158 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_159 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'h9f == io_addrb) begin // @[RAM.scala 50:23]
        mem_159 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_160 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha0 == io_addrb) begin // @[RAM.scala 50:23]
        mem_160 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_161 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha1 == io_addrb) begin // @[RAM.scala 50:23]
        mem_161 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_162 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha2 == io_addrb) begin // @[RAM.scala 50:23]
        mem_162 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_163 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha3 == io_addrb) begin // @[RAM.scala 50:23]
        mem_163 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_164 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha4 == io_addrb) begin // @[RAM.scala 50:23]
        mem_164 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_165 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha5 == io_addrb) begin // @[RAM.scala 50:23]
        mem_165 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_166 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha6 == io_addrb) begin // @[RAM.scala 50:23]
        mem_166 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_167 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha7 == io_addrb) begin // @[RAM.scala 50:23]
        mem_167 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_168 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha8 == io_addrb) begin // @[RAM.scala 50:23]
        mem_168 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_169 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'ha9 == io_addrb) begin // @[RAM.scala 50:23]
        mem_169 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_170 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'haa == io_addrb) begin // @[RAM.scala 50:23]
        mem_170 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_171 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hab == io_addrb) begin // @[RAM.scala 50:23]
        mem_171 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_172 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hac == io_addrb) begin // @[RAM.scala 50:23]
        mem_172 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_173 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'had == io_addrb) begin // @[RAM.scala 50:23]
        mem_173 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_174 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hae == io_addrb) begin // @[RAM.scala 50:23]
        mem_174 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_175 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'haf == io_addrb) begin // @[RAM.scala 50:23]
        mem_175 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_176 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb0 == io_addrb) begin // @[RAM.scala 50:23]
        mem_176 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_177 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb1 == io_addrb) begin // @[RAM.scala 50:23]
        mem_177 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_178 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb2 == io_addrb) begin // @[RAM.scala 50:23]
        mem_178 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_179 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb3 == io_addrb) begin // @[RAM.scala 50:23]
        mem_179 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_180 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb4 == io_addrb) begin // @[RAM.scala 50:23]
        mem_180 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_181 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb5 == io_addrb) begin // @[RAM.scala 50:23]
        mem_181 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_182 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb6 == io_addrb) begin // @[RAM.scala 50:23]
        mem_182 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_183 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb7 == io_addrb) begin // @[RAM.scala 50:23]
        mem_183 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_184 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb8 == io_addrb) begin // @[RAM.scala 50:23]
        mem_184 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_185 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hb9 == io_addrb) begin // @[RAM.scala 50:23]
        mem_185 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_186 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hba == io_addrb) begin // @[RAM.scala 50:23]
        mem_186 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_187 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hbb == io_addrb) begin // @[RAM.scala 50:23]
        mem_187 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_188 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hbc == io_addrb) begin // @[RAM.scala 50:23]
        mem_188 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_189 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hbd == io_addrb) begin // @[RAM.scala 50:23]
        mem_189 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_190 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hbe == io_addrb) begin // @[RAM.scala 50:23]
        mem_190 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_191 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hbf == io_addrb) begin // @[RAM.scala 50:23]
        mem_191 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_192 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc0 == io_addrb) begin // @[RAM.scala 50:23]
        mem_192 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_193 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc1 == io_addrb) begin // @[RAM.scala 50:23]
        mem_193 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_194 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc2 == io_addrb) begin // @[RAM.scala 50:23]
        mem_194 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_195 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc3 == io_addrb) begin // @[RAM.scala 50:23]
        mem_195 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_196 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc4 == io_addrb) begin // @[RAM.scala 50:23]
        mem_196 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_197 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc5 == io_addrb) begin // @[RAM.scala 50:23]
        mem_197 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_198 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc6 == io_addrb) begin // @[RAM.scala 50:23]
        mem_198 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_199 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc7 == io_addrb) begin // @[RAM.scala 50:23]
        mem_199 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_200 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc8 == io_addrb) begin // @[RAM.scala 50:23]
        mem_200 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_201 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hc9 == io_addrb) begin // @[RAM.scala 50:23]
        mem_201 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_202 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hca == io_addrb) begin // @[RAM.scala 50:23]
        mem_202 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_203 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hcb == io_addrb) begin // @[RAM.scala 50:23]
        mem_203 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_204 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hcc == io_addrb) begin // @[RAM.scala 50:23]
        mem_204 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_205 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hcd == io_addrb) begin // @[RAM.scala 50:23]
        mem_205 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_206 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hce == io_addrb) begin // @[RAM.scala 50:23]
        mem_206 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_207 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hcf == io_addrb) begin // @[RAM.scala 50:23]
        mem_207 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_208 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd0 == io_addrb) begin // @[RAM.scala 50:23]
        mem_208 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_209 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd1 == io_addrb) begin // @[RAM.scala 50:23]
        mem_209 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_210 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd2 == io_addrb) begin // @[RAM.scala 50:23]
        mem_210 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_211 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd3 == io_addrb) begin // @[RAM.scala 50:23]
        mem_211 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_212 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd4 == io_addrb) begin // @[RAM.scala 50:23]
        mem_212 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_213 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd5 == io_addrb) begin // @[RAM.scala 50:23]
        mem_213 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_214 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd6 == io_addrb) begin // @[RAM.scala 50:23]
        mem_214 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_215 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd7 == io_addrb) begin // @[RAM.scala 50:23]
        mem_215 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_216 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd8 == io_addrb) begin // @[RAM.scala 50:23]
        mem_216 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_217 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hd9 == io_addrb) begin // @[RAM.scala 50:23]
        mem_217 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_218 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hda == io_addrb) begin // @[RAM.scala 50:23]
        mem_218 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_219 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hdb == io_addrb) begin // @[RAM.scala 50:23]
        mem_219 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_220 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hdc == io_addrb) begin // @[RAM.scala 50:23]
        mem_220 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_221 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hdd == io_addrb) begin // @[RAM.scala 50:23]
        mem_221 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_222 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hde == io_addrb) begin // @[RAM.scala 50:23]
        mem_222 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_223 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hdf == io_addrb) begin // @[RAM.scala 50:23]
        mem_223 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_224 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he0 == io_addrb) begin // @[RAM.scala 50:23]
        mem_224 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_225 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he1 == io_addrb) begin // @[RAM.scala 50:23]
        mem_225 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_226 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he2 == io_addrb) begin // @[RAM.scala 50:23]
        mem_226 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_227 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he3 == io_addrb) begin // @[RAM.scala 50:23]
        mem_227 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_228 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he4 == io_addrb) begin // @[RAM.scala 50:23]
        mem_228 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_229 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he5 == io_addrb) begin // @[RAM.scala 50:23]
        mem_229 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_230 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he6 == io_addrb) begin // @[RAM.scala 50:23]
        mem_230 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_231 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he7 == io_addrb) begin // @[RAM.scala 50:23]
        mem_231 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_232 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he8 == io_addrb) begin // @[RAM.scala 50:23]
        mem_232 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_233 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'he9 == io_addrb) begin // @[RAM.scala 50:23]
        mem_233 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_234 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hea == io_addrb) begin // @[RAM.scala 50:23]
        mem_234 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_235 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'heb == io_addrb) begin // @[RAM.scala 50:23]
        mem_235 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_236 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hec == io_addrb) begin // @[RAM.scala 50:23]
        mem_236 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_237 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hed == io_addrb) begin // @[RAM.scala 50:23]
        mem_237 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_238 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hee == io_addrb) begin // @[RAM.scala 50:23]
        mem_238 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_239 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hef == io_addrb) begin // @[RAM.scala 50:23]
        mem_239 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_240 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf0 == io_addrb) begin // @[RAM.scala 50:23]
        mem_240 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_241 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf1 == io_addrb) begin // @[RAM.scala 50:23]
        mem_241 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_242 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf2 == io_addrb) begin // @[RAM.scala 50:23]
        mem_242 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_243 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf3 == io_addrb) begin // @[RAM.scala 50:23]
        mem_243 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_244 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf4 == io_addrb) begin // @[RAM.scala 50:23]
        mem_244 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_245 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf5 == io_addrb) begin // @[RAM.scala 50:23]
        mem_245 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_246 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf6 == io_addrb) begin // @[RAM.scala 50:23]
        mem_246 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_247 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf7 == io_addrb) begin // @[RAM.scala 50:23]
        mem_247 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_248 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf8 == io_addrb) begin // @[RAM.scala 50:23]
        mem_248 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_249 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hf9 == io_addrb) begin // @[RAM.scala 50:23]
        mem_249 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_250 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hfa == io_addrb) begin // @[RAM.scala 50:23]
        mem_250 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_251 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hfb == io_addrb) begin // @[RAM.scala 50:23]
        mem_251 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_252 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hfc == io_addrb) begin // @[RAM.scala 50:23]
        mem_252 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_253 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hfd == io_addrb) begin // @[RAM.scala 50:23]
        mem_253 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_254 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hfe == io_addrb) begin // @[RAM.scala 50:23]
        mem_254 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (reset) begin // @[RAM.scala 41:22]
      mem_255 <= 22'h0; // @[RAM.scala 41:22]
    end else if (io_web) begin // @[RAM.scala 49:18]
      if (8'hff == io_addrb) begin // @[RAM.scala 50:23]
        mem_255 <= io_dinb; // @[RAM.scala 50:23]
      end
    end
    if (8'hff == io_addra) begin // @[RAM.scala 43:24]
      io_douta_REG <= mem_255; // @[RAM.scala 43:24]
    end else if (8'hfe == io_addra) begin // @[RAM.scala 43:24]
      io_douta_REG <= mem_254; // @[RAM.scala 43:24]
    end else if (8'hfd == io_addra) begin // @[RAM.scala 43:24]
      io_douta_REG <= mem_253; // @[RAM.scala 43:24]
    end else if (8'hfc == io_addra) begin // @[RAM.scala 43:24]
      io_douta_REG <= mem_252; // @[RAM.scala 43:24]
    end else begin
      io_douta_REG <= _GEN_251;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0 = _RAND_0[21:0];
  _RAND_1 = {1{`RANDOM}};
  mem_1 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  mem_2 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  mem_3 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  mem_4 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  mem_5 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  mem_6 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  mem_7 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  mem_8 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  mem_9 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  mem_10 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  mem_11 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  mem_12 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  mem_13 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  mem_14 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  mem_15 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  mem_16 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  mem_17 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  mem_18 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  mem_19 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  mem_20 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  mem_21 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  mem_22 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  mem_23 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  mem_24 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  mem_25 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  mem_26 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  mem_27 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  mem_28 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  mem_29 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  mem_30 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  mem_31 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  mem_32 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  mem_33 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  mem_34 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  mem_35 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  mem_36 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  mem_37 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  mem_38 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  mem_39 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  mem_40 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  mem_41 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  mem_42 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  mem_43 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  mem_44 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  mem_45 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  mem_46 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  mem_47 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  mem_48 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  mem_49 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  mem_50 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  mem_51 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  mem_52 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  mem_53 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  mem_54 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  mem_55 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  mem_56 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  mem_57 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  mem_58 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  mem_59 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  mem_60 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  mem_61 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  mem_62 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  mem_63 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  mem_64 = _RAND_64[21:0];
  _RAND_65 = {1{`RANDOM}};
  mem_65 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  mem_66 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  mem_67 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  mem_68 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  mem_69 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  mem_70 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  mem_71 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  mem_72 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  mem_73 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  mem_74 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  mem_75 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  mem_76 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  mem_77 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  mem_78 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  mem_79 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  mem_80 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  mem_81 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  mem_82 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  mem_83 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  mem_84 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  mem_85 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  mem_86 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  mem_87 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  mem_88 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  mem_89 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  mem_90 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  mem_91 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  mem_92 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  mem_93 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  mem_94 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  mem_95 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  mem_96 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  mem_97 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  mem_98 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  mem_99 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  mem_100 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  mem_101 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  mem_102 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  mem_103 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  mem_104 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  mem_105 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  mem_106 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  mem_107 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  mem_108 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  mem_109 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  mem_110 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  mem_111 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  mem_112 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  mem_113 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  mem_114 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  mem_115 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  mem_116 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  mem_117 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  mem_118 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  mem_119 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  mem_120 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  mem_121 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  mem_122 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  mem_123 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  mem_124 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  mem_125 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  mem_126 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  mem_127 = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  mem_128 = _RAND_128[21:0];
  _RAND_129 = {1{`RANDOM}};
  mem_129 = _RAND_129[21:0];
  _RAND_130 = {1{`RANDOM}};
  mem_130 = _RAND_130[21:0];
  _RAND_131 = {1{`RANDOM}};
  mem_131 = _RAND_131[21:0];
  _RAND_132 = {1{`RANDOM}};
  mem_132 = _RAND_132[21:0];
  _RAND_133 = {1{`RANDOM}};
  mem_133 = _RAND_133[21:0];
  _RAND_134 = {1{`RANDOM}};
  mem_134 = _RAND_134[21:0];
  _RAND_135 = {1{`RANDOM}};
  mem_135 = _RAND_135[21:0];
  _RAND_136 = {1{`RANDOM}};
  mem_136 = _RAND_136[21:0];
  _RAND_137 = {1{`RANDOM}};
  mem_137 = _RAND_137[21:0];
  _RAND_138 = {1{`RANDOM}};
  mem_138 = _RAND_138[21:0];
  _RAND_139 = {1{`RANDOM}};
  mem_139 = _RAND_139[21:0];
  _RAND_140 = {1{`RANDOM}};
  mem_140 = _RAND_140[21:0];
  _RAND_141 = {1{`RANDOM}};
  mem_141 = _RAND_141[21:0];
  _RAND_142 = {1{`RANDOM}};
  mem_142 = _RAND_142[21:0];
  _RAND_143 = {1{`RANDOM}};
  mem_143 = _RAND_143[21:0];
  _RAND_144 = {1{`RANDOM}};
  mem_144 = _RAND_144[21:0];
  _RAND_145 = {1{`RANDOM}};
  mem_145 = _RAND_145[21:0];
  _RAND_146 = {1{`RANDOM}};
  mem_146 = _RAND_146[21:0];
  _RAND_147 = {1{`RANDOM}};
  mem_147 = _RAND_147[21:0];
  _RAND_148 = {1{`RANDOM}};
  mem_148 = _RAND_148[21:0];
  _RAND_149 = {1{`RANDOM}};
  mem_149 = _RAND_149[21:0];
  _RAND_150 = {1{`RANDOM}};
  mem_150 = _RAND_150[21:0];
  _RAND_151 = {1{`RANDOM}};
  mem_151 = _RAND_151[21:0];
  _RAND_152 = {1{`RANDOM}};
  mem_152 = _RAND_152[21:0];
  _RAND_153 = {1{`RANDOM}};
  mem_153 = _RAND_153[21:0];
  _RAND_154 = {1{`RANDOM}};
  mem_154 = _RAND_154[21:0];
  _RAND_155 = {1{`RANDOM}};
  mem_155 = _RAND_155[21:0];
  _RAND_156 = {1{`RANDOM}};
  mem_156 = _RAND_156[21:0];
  _RAND_157 = {1{`RANDOM}};
  mem_157 = _RAND_157[21:0];
  _RAND_158 = {1{`RANDOM}};
  mem_158 = _RAND_158[21:0];
  _RAND_159 = {1{`RANDOM}};
  mem_159 = _RAND_159[21:0];
  _RAND_160 = {1{`RANDOM}};
  mem_160 = _RAND_160[21:0];
  _RAND_161 = {1{`RANDOM}};
  mem_161 = _RAND_161[21:0];
  _RAND_162 = {1{`RANDOM}};
  mem_162 = _RAND_162[21:0];
  _RAND_163 = {1{`RANDOM}};
  mem_163 = _RAND_163[21:0];
  _RAND_164 = {1{`RANDOM}};
  mem_164 = _RAND_164[21:0];
  _RAND_165 = {1{`RANDOM}};
  mem_165 = _RAND_165[21:0];
  _RAND_166 = {1{`RANDOM}};
  mem_166 = _RAND_166[21:0];
  _RAND_167 = {1{`RANDOM}};
  mem_167 = _RAND_167[21:0];
  _RAND_168 = {1{`RANDOM}};
  mem_168 = _RAND_168[21:0];
  _RAND_169 = {1{`RANDOM}};
  mem_169 = _RAND_169[21:0];
  _RAND_170 = {1{`RANDOM}};
  mem_170 = _RAND_170[21:0];
  _RAND_171 = {1{`RANDOM}};
  mem_171 = _RAND_171[21:0];
  _RAND_172 = {1{`RANDOM}};
  mem_172 = _RAND_172[21:0];
  _RAND_173 = {1{`RANDOM}};
  mem_173 = _RAND_173[21:0];
  _RAND_174 = {1{`RANDOM}};
  mem_174 = _RAND_174[21:0];
  _RAND_175 = {1{`RANDOM}};
  mem_175 = _RAND_175[21:0];
  _RAND_176 = {1{`RANDOM}};
  mem_176 = _RAND_176[21:0];
  _RAND_177 = {1{`RANDOM}};
  mem_177 = _RAND_177[21:0];
  _RAND_178 = {1{`RANDOM}};
  mem_178 = _RAND_178[21:0];
  _RAND_179 = {1{`RANDOM}};
  mem_179 = _RAND_179[21:0];
  _RAND_180 = {1{`RANDOM}};
  mem_180 = _RAND_180[21:0];
  _RAND_181 = {1{`RANDOM}};
  mem_181 = _RAND_181[21:0];
  _RAND_182 = {1{`RANDOM}};
  mem_182 = _RAND_182[21:0];
  _RAND_183 = {1{`RANDOM}};
  mem_183 = _RAND_183[21:0];
  _RAND_184 = {1{`RANDOM}};
  mem_184 = _RAND_184[21:0];
  _RAND_185 = {1{`RANDOM}};
  mem_185 = _RAND_185[21:0];
  _RAND_186 = {1{`RANDOM}};
  mem_186 = _RAND_186[21:0];
  _RAND_187 = {1{`RANDOM}};
  mem_187 = _RAND_187[21:0];
  _RAND_188 = {1{`RANDOM}};
  mem_188 = _RAND_188[21:0];
  _RAND_189 = {1{`RANDOM}};
  mem_189 = _RAND_189[21:0];
  _RAND_190 = {1{`RANDOM}};
  mem_190 = _RAND_190[21:0];
  _RAND_191 = {1{`RANDOM}};
  mem_191 = _RAND_191[21:0];
  _RAND_192 = {1{`RANDOM}};
  mem_192 = _RAND_192[21:0];
  _RAND_193 = {1{`RANDOM}};
  mem_193 = _RAND_193[21:0];
  _RAND_194 = {1{`RANDOM}};
  mem_194 = _RAND_194[21:0];
  _RAND_195 = {1{`RANDOM}};
  mem_195 = _RAND_195[21:0];
  _RAND_196 = {1{`RANDOM}};
  mem_196 = _RAND_196[21:0];
  _RAND_197 = {1{`RANDOM}};
  mem_197 = _RAND_197[21:0];
  _RAND_198 = {1{`RANDOM}};
  mem_198 = _RAND_198[21:0];
  _RAND_199 = {1{`RANDOM}};
  mem_199 = _RAND_199[21:0];
  _RAND_200 = {1{`RANDOM}};
  mem_200 = _RAND_200[21:0];
  _RAND_201 = {1{`RANDOM}};
  mem_201 = _RAND_201[21:0];
  _RAND_202 = {1{`RANDOM}};
  mem_202 = _RAND_202[21:0];
  _RAND_203 = {1{`RANDOM}};
  mem_203 = _RAND_203[21:0];
  _RAND_204 = {1{`RANDOM}};
  mem_204 = _RAND_204[21:0];
  _RAND_205 = {1{`RANDOM}};
  mem_205 = _RAND_205[21:0];
  _RAND_206 = {1{`RANDOM}};
  mem_206 = _RAND_206[21:0];
  _RAND_207 = {1{`RANDOM}};
  mem_207 = _RAND_207[21:0];
  _RAND_208 = {1{`RANDOM}};
  mem_208 = _RAND_208[21:0];
  _RAND_209 = {1{`RANDOM}};
  mem_209 = _RAND_209[21:0];
  _RAND_210 = {1{`RANDOM}};
  mem_210 = _RAND_210[21:0];
  _RAND_211 = {1{`RANDOM}};
  mem_211 = _RAND_211[21:0];
  _RAND_212 = {1{`RANDOM}};
  mem_212 = _RAND_212[21:0];
  _RAND_213 = {1{`RANDOM}};
  mem_213 = _RAND_213[21:0];
  _RAND_214 = {1{`RANDOM}};
  mem_214 = _RAND_214[21:0];
  _RAND_215 = {1{`RANDOM}};
  mem_215 = _RAND_215[21:0];
  _RAND_216 = {1{`RANDOM}};
  mem_216 = _RAND_216[21:0];
  _RAND_217 = {1{`RANDOM}};
  mem_217 = _RAND_217[21:0];
  _RAND_218 = {1{`RANDOM}};
  mem_218 = _RAND_218[21:0];
  _RAND_219 = {1{`RANDOM}};
  mem_219 = _RAND_219[21:0];
  _RAND_220 = {1{`RANDOM}};
  mem_220 = _RAND_220[21:0];
  _RAND_221 = {1{`RANDOM}};
  mem_221 = _RAND_221[21:0];
  _RAND_222 = {1{`RANDOM}};
  mem_222 = _RAND_222[21:0];
  _RAND_223 = {1{`RANDOM}};
  mem_223 = _RAND_223[21:0];
  _RAND_224 = {1{`RANDOM}};
  mem_224 = _RAND_224[21:0];
  _RAND_225 = {1{`RANDOM}};
  mem_225 = _RAND_225[21:0];
  _RAND_226 = {1{`RANDOM}};
  mem_226 = _RAND_226[21:0];
  _RAND_227 = {1{`RANDOM}};
  mem_227 = _RAND_227[21:0];
  _RAND_228 = {1{`RANDOM}};
  mem_228 = _RAND_228[21:0];
  _RAND_229 = {1{`RANDOM}};
  mem_229 = _RAND_229[21:0];
  _RAND_230 = {1{`RANDOM}};
  mem_230 = _RAND_230[21:0];
  _RAND_231 = {1{`RANDOM}};
  mem_231 = _RAND_231[21:0];
  _RAND_232 = {1{`RANDOM}};
  mem_232 = _RAND_232[21:0];
  _RAND_233 = {1{`RANDOM}};
  mem_233 = _RAND_233[21:0];
  _RAND_234 = {1{`RANDOM}};
  mem_234 = _RAND_234[21:0];
  _RAND_235 = {1{`RANDOM}};
  mem_235 = _RAND_235[21:0];
  _RAND_236 = {1{`RANDOM}};
  mem_236 = _RAND_236[21:0];
  _RAND_237 = {1{`RANDOM}};
  mem_237 = _RAND_237[21:0];
  _RAND_238 = {1{`RANDOM}};
  mem_238 = _RAND_238[21:0];
  _RAND_239 = {1{`RANDOM}};
  mem_239 = _RAND_239[21:0];
  _RAND_240 = {1{`RANDOM}};
  mem_240 = _RAND_240[21:0];
  _RAND_241 = {1{`RANDOM}};
  mem_241 = _RAND_241[21:0];
  _RAND_242 = {1{`RANDOM}};
  mem_242 = _RAND_242[21:0];
  _RAND_243 = {1{`RANDOM}};
  mem_243 = _RAND_243[21:0];
  _RAND_244 = {1{`RANDOM}};
  mem_244 = _RAND_244[21:0];
  _RAND_245 = {1{`RANDOM}};
  mem_245 = _RAND_245[21:0];
  _RAND_246 = {1{`RANDOM}};
  mem_246 = _RAND_246[21:0];
  _RAND_247 = {1{`RANDOM}};
  mem_247 = _RAND_247[21:0];
  _RAND_248 = {1{`RANDOM}};
  mem_248 = _RAND_248[21:0];
  _RAND_249 = {1{`RANDOM}};
  mem_249 = _RAND_249[21:0];
  _RAND_250 = {1{`RANDOM}};
  mem_250 = _RAND_250[21:0];
  _RAND_251 = {1{`RANDOM}};
  mem_251 = _RAND_251[21:0];
  _RAND_252 = {1{`RANDOM}};
  mem_252 = _RAND_252[21:0];
  _RAND_253 = {1{`RANDOM}};
  mem_253 = _RAND_253[21:0];
  _RAND_254 = {1{`RANDOM}};
  mem_254 = _RAND_254[21:0];
  _RAND_255 = {1{`RANDOM}};
  mem_255 = _RAND_255[21:0];
  _RAND_256 = {1{`RANDOM}};
  io_douta_REG = _RAND_256[21:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DualPortBRAM_2(
  input         clock,
  input         reset,
  input         io_web,
  input  [7:0]  io_addra,
  input  [7:0]  io_addrb,
  input  [21:0] io_dinb,
  output [21:0] io_douta
);
  wire  sim_dual_port_bram_clock; // @[RAM.scala 30:40]
  wire  sim_dual_port_bram_reset; // @[RAM.scala 30:40]
  wire  sim_dual_port_bram_io_web; // @[RAM.scala 30:40]
  wire [7:0] sim_dual_port_bram_io_addra; // @[RAM.scala 30:40]
  wire [7:0] sim_dual_port_bram_io_addrb; // @[RAM.scala 30:40]
  wire [21:0] sim_dual_port_bram_io_dinb; // @[RAM.scala 30:40]
  wire [21:0] sim_dual_port_bram_io_douta; // @[RAM.scala 30:40]
  SimDualPortBRAM_2 sim_dual_port_bram ( // @[RAM.scala 30:40]
    .clock(sim_dual_port_bram_clock),
    .reset(sim_dual_port_bram_reset),
    .io_web(sim_dual_port_bram_io_web),
    .io_addra(sim_dual_port_bram_io_addra),
    .io_addrb(sim_dual_port_bram_io_addrb),
    .io_dinb(sim_dual_port_bram_io_dinb),
    .io_douta(sim_dual_port_bram_io_douta)
  );
  assign io_douta = sim_dual_port_bram_io_douta; // @[RAM.scala 31:31]
  assign sim_dual_port_bram_clock = clock;
  assign sim_dual_port_bram_reset = reset;
  assign sim_dual_port_bram_io_web = io_web; // @[RAM.scala 31:31]
  assign sim_dual_port_bram_io_addra = io_addra; // @[RAM.scala 31:31]
  assign sim_dual_port_bram_io_addrb = io_addrb; // @[RAM.scala 31:31]
  assign sim_dual_port_bram_io_dinb = io_dinb; // @[RAM.scala 31:31]
endmodule
module MetaDataBRAM(
  input         clock,
  input         reset,
  input  [7:0]  io_indexFetch,
  input  [7:0]  io_indexUpdate,
  input  [19:0] io_tagUpdate,
  input         io_update,
  input         io_write,
  output        io_hit,
  output [19:0] io_tagFetch
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  blk_clock; // @[DCache.scala 28:19]
  wire  blk_reset; // @[DCache.scala 28:19]
  wire  blk_io_web; // @[DCache.scala 28:19]
  wire [7:0] blk_io_addra; // @[DCache.scala 28:19]
  wire [7:0] blk_io_addrb; // @[DCache.scala 28:19]
  wire [21:0] blk_io_dinb; // @[DCache.scala 28:19]
  wire [21:0] blk_io_douta; // @[DCache.scala 28:19]
  reg  dout_REG; // @[DCache.scala 31:25]
  reg [21:0] dout_REG_1; // @[DCache.scala 31:79]
  wire [21:0] dout = dout_REG ? dout_REG_1 : blk_io_douta; // @[DCache.scala 31:17]
  wire  v = dout[20]; // @[DCache.scala 32:15]
  wire [19:0] tag = dout[19:0]; // @[DCache.scala 33:17]
  wire [1:0] blk_io_dinb_hi = {io_write,1'h1}; // @[Cat.scala 30:58]
  DualPortBRAM_2 blk ( // @[DCache.scala 28:19]
    .clock(blk_clock),
    .reset(blk_reset),
    .io_web(blk_io_web),
    .io_addra(blk_io_addra),
    .io_addrb(blk_io_addrb),
    .io_dinb(blk_io_dinb),
    .io_douta(blk_io_douta)
  );
  assign io_hit = v & io_tagUpdate == tag; // @[DCache.scala 47:21]
  assign io_tagFetch = dout[19:0]; // @[DCache.scala 33:17]
  assign blk_clock = clock;
  assign blk_reset = reset;
  assign blk_io_web = io_update; // @[DCache.scala 42:16]
  assign blk_io_addra = io_indexFetch; // @[DCache.scala 39:16]
  assign blk_io_addrb = io_indexUpdate; // @[DCache.scala 43:16]
  assign blk_io_dinb = {blk_io_dinb_hi,io_tagUpdate}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    dout_REG <= blk_io_web & blk_io_addra == blk_io_addrb; // @[DCache.scala 31:37]
    dout_REG_1 <= blk_io_dinb; // @[DCache.scala 31:79]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dout_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  dout_REG_1 = _RAND_1[21:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCache(
  input          clock,
  input          reset,
  output         io_cpu_req_ready,
  input          io_cpu_req_valid,
  input  [31:0]  io_cpu_req_bits_addr,
  input          io_cpu_req_bits_wen,
  input  [31:0]  io_cpu_req_bits_wdata,
  input  [1:0]   io_cpu_req_bits_mtype,
  output         io_cpu_resp_valid,
  output [31:0]  io_cpu_resp_bits_rdata,
  output [31:0]  io_bar_req_bits_addr,
  output         io_bar_req_bits_wen,
  output [127:0] io_bar_req_bits_wdata,
  output [1:0]   io_bar_req_bits_mtype,
  input  [127:0] io_bar_resp_bits_rdata,
  output         io_dbg_hit,
  output         io_dbg_hitWay,
  output         io_dbg_replaceWay
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  wire  data_0_clock; // @[DCache.scala 54:48]
  wire  data_0_reset; // @[DCache.scala 54:48]
  wire  data_0_io_web; // @[DCache.scala 54:48]
  wire [7:0] data_0_io_addra; // @[DCache.scala 54:48]
  wire [7:0] data_0_io_addrb; // @[DCache.scala 54:48]
  wire [127:0] data_0_io_dinb; // @[DCache.scala 54:48]
  wire [127:0] data_0_io_douta; // @[DCache.scala 54:48]
  wire  data_1_clock; // @[DCache.scala 54:48]
  wire  data_1_reset; // @[DCache.scala 54:48]
  wire  data_1_io_web; // @[DCache.scala 54:48]
  wire [7:0] data_1_io_addra; // @[DCache.scala 54:48]
  wire [7:0] data_1_io_addrb; // @[DCache.scala 54:48]
  wire [127:0] data_1_io_dinb; // @[DCache.scala 54:48]
  wire [127:0] data_1_io_douta; // @[DCache.scala 54:48]
  wire  meta_0_clock; // @[DCache.scala 55:48]
  wire  meta_0_reset; // @[DCache.scala 55:48]
  wire [7:0] meta_0_io_indexFetch; // @[DCache.scala 55:48]
  wire [7:0] meta_0_io_indexUpdate; // @[DCache.scala 55:48]
  wire [19:0] meta_0_io_tagUpdate; // @[DCache.scala 55:48]
  wire  meta_0_io_update; // @[DCache.scala 55:48]
  wire  meta_0_io_write; // @[DCache.scala 55:48]
  wire  meta_0_io_hit; // @[DCache.scala 55:48]
  wire [19:0] meta_0_io_tagFetch; // @[DCache.scala 55:48]
  wire  meta_1_clock; // @[DCache.scala 55:48]
  wire  meta_1_reset; // @[DCache.scala 55:48]
  wire [7:0] meta_1_io_indexFetch; // @[DCache.scala 55:48]
  wire [7:0] meta_1_io_indexUpdate; // @[DCache.scala 55:48]
  wire [19:0] meta_1_io_tagUpdate; // @[DCache.scala 55:48]
  wire  meta_1_io_update; // @[DCache.scala 55:48]
  wire  meta_1_io_write; // @[DCache.scala 55:48]
  wire  meta_1_io_hit; // @[DCache.scala 55:48]
  wire [19:0] meta_1_io_tagFetch; // @[DCache.scala 55:48]
  wire [1:0] arOffset = io_cpu_req_bits_addr[3:2]; // @[DCache.scala 64:40]
  wire [7:0] arIndex = io_cpu_req_bits_addr[11:4]; // @[DCache.scala 65:40]
  wire [19:0] arTag = io_cpu_req_bits_addr[31:12]; // @[DCache.scala 66:40]
  reg  mpValid; // @[DCache.scala 85:26]
  reg  mpState; // @[DCache.scala 163:26]
  wire  _T_31 = ~mpState; // @[Conditional.scala 37:30]
  wire  mpWriteCache = mpValid & mpState; // @[DCache.scala 165:29]
  wire  _GEN_57 = mpState & mpWriteCache; // @[Conditional.scala 39:67 DCache.scala 207:29 DCache.scala 195:17]
  wire  _GEN_61 = _T_31 ? 1'h0 : _GEN_57; // @[Conditional.scala 40:58 DCache.scala 195:17]
  wire  mpRespValid = mpValid & _GEN_61; // @[DCache.scala 196:20 DCache.scala 195:17]
  wire  mpStall = mpValid & ~mpRespValid; // @[DCache.scala 87:27]
  wire  _hpReq_T = ~mpStall; // @[DCache.scala 75:50]
  reg [31:0] hpReq_addr; // @[Reg.scala 15:16]
  reg  hpReq_wen; // @[Reg.scala 15:16]
  reg [31:0] hpReq_wdata; // @[Reg.scala 15:16]
  reg [1:0] hpReq_mtype; // @[Reg.scala 15:16]
  reg [7:0] hpIndex; // @[Reg.scala 15:16]
  reg [19:0] hpTag; // @[Reg.scala 15:16]
  reg [1:0] hpOffset; // @[Reg.scala 15:16]
  reg  hpValid; // @[DCache.scala 79:30]
  wire  _hpRespValid_T = meta_0_io_hit | meta_1_io_hit; // @[DCache.scala 80:50]
  wire  hpRespValid = hpValid & (meta_0_io_hit | meta_1_io_hit); // @[DCache.scala 80:31]
  reg  mpReq_wen; // @[DCache.scala 83:26]
  reg [31:0] mpReq_wdata; // @[DCache.scala 83:26]
  reg [31:0] mpDirtyAddr; // @[DCache.scala 91:27]
  reg [127:0] mpDirtyData; // @[DCache.scala 92:27]
  reg [3:0] mpOffset; // @[DCache.scala 93:27]
  reg [7:0] mpIndex; // @[DCache.scala 94:27]
  reg [19:0] mpTag; // @[DCache.scala 95:27]
  wire [31:0] mpRefillAddr = {mpTag,mpIndex,4'h0}; // @[Cat.scala 30:58]
  reg [31:0] mpMask; // @[DCache.scala 97:23]
  reg [4:0] mpShift; // @[DCache.scala 98:23]
  wire  _hpValid_T_1 = hpValid & ~_hpRespValid_T; // @[DCache.scala 111:29]
  reg  REG; // @[DCache.scala 118:38]
  wire [127:0] _WIRE_1 = data_0_io_dinb;
  reg [31:0] REG_1_0; // @[DCache.scala 119:40]
  reg [31:0] REG_1_1; // @[DCache.scala 119:40]
  reg [31:0] REG_1_2; // @[DCache.scala 119:40]
  reg [31:0] REG_1_3; // @[DCache.scala 119:40]
  wire [127:0] _WIRE_3 = data_0_io_douta;
  wire [31:0] hpFetchLine_0_0 = REG ? REG_1_0 : _WIRE_3[31:0]; // @[DCache.scala 118:30]
  wire [31:0] hpFetchLine_0_1 = REG ? REG_1_1 : _WIRE_3[63:32]; // @[DCache.scala 118:30]
  wire [31:0] hpFetchLine_0_2 = REG ? REG_1_2 : _WIRE_3[95:64]; // @[DCache.scala 118:30]
  wire [31:0] hpFetchLine_0_3 = REG ? REG_1_3 : _WIRE_3[127:96]; // @[DCache.scala 118:30]
  reg  REG_2; // @[DCache.scala 118:38]
  wire [127:0] _WIRE_5 = data_1_io_dinb;
  reg [31:0] REG_3_0; // @[DCache.scala 119:40]
  reg [31:0] REG_3_1; // @[DCache.scala 119:40]
  reg [31:0] REG_3_2; // @[DCache.scala 119:40]
  reg [31:0] REG_3_3; // @[DCache.scala 119:40]
  wire [127:0] _WIRE_7 = data_1_io_douta;
  wire [31:0] hpFetchLine_1_0 = REG_2 ? REG_3_0 : _WIRE_7[31:0]; // @[DCache.scala 118:30]
  wire [31:0] hpFetchLine_1_1 = REG_2 ? REG_3_1 : _WIRE_7[63:32]; // @[DCache.scala 118:30]
  wire [31:0] hpFetchLine_1_2 = REG_2 ? REG_3_2 : _WIRE_7[95:64]; // @[DCache.scala 118:30]
  wire [31:0] hpFetchLine_1_3 = REG_2 ? REG_3_3 : _WIRE_7[127:96]; // @[DCache.scala 118:30]
  wire [31:0] _hpMask_T_1 = 2'h0 == hpReq_mtype ? 32'hff : 32'hffffffff; // @[Mux.scala 80:57]
  wire [31:0] hpMask = 2'h1 == hpReq_mtype ? 32'hffff : _hpMask_T_1; // @[Mux.scala 80:57]
  wire [4:0] hpShift = {hpReq_addr[1:0], 3'h0}; // @[DCache.scala 129:50]
  wire [31:0] _hpWriteWord_0_T = hpMask & hpReq_wdata; // @[DCache.scala 135:36]
  wire [62:0] _GEN_66 = {{31'd0}, _hpWriteWord_0_T}; // @[DCache.scala 135:51]
  wire [62:0] _hpWriteWord_0_T_1 = _GEN_66 << hpShift; // @[DCache.scala 135:51]
  wire [62:0] _GEN_67 = {{31'd0}, hpMask}; // @[DCache.scala 135:85]
  wire [62:0] _hpWriteWord_0_T_2 = _GEN_67 << hpShift; // @[DCache.scala 135:85]
  wire [62:0] _hpWriteWord_0_T_3 = ~_hpWriteWord_0_T_2; // @[DCache.scala 135:76]
  wire [31:0] _GEN_8 = 2'h1 == hpOffset ? hpFetchLine_0_1 : hpFetchLine_0_0; // @[DCache.scala 135:107 DCache.scala 135:107]
  wire [31:0] _GEN_9 = 2'h2 == hpOffset ? hpFetchLine_0_2 : _GEN_8; // @[DCache.scala 135:107 DCache.scala 135:107]
  wire [31:0] _GEN_10 = 2'h3 == hpOffset ? hpFetchLine_0_3 : _GEN_9; // @[DCache.scala 135:107 DCache.scala 135:107]
  wire [62:0] _GEN_68 = {{31'd0}, _GEN_10}; // @[DCache.scala 135:107]
  wire [62:0] _hpWriteWord_0_T_4 = _hpWriteWord_0_T_3 & _GEN_68; // @[DCache.scala 135:107]
  wire [62:0] _hpWriteWord_0_T_5 = _hpWriteWord_0_T_1 | _hpWriteWord_0_T_4; // @[DCache.scala 135:72]
  wire [31:0] hpWriteWord_0 = _hpWriteWord_0_T_5[31:0]; // @[DCache.scala 130:27 DCache.scala 135:24]
  wire [31:0] hpWriteLine_0_0 = 2'h0 == hpOffset ? hpWriteWord_0 : hpFetchLine_0_0; // @[DCache.scala 138:34 DCache.scala 138:34 DCache.scala 137:24]
  wire [31:0] hpWriteLine_0_1 = 2'h1 == hpOffset ? hpWriteWord_0 : hpFetchLine_0_1; // @[DCache.scala 138:34 DCache.scala 138:34 DCache.scala 137:24]
  wire [31:0] hpWriteLine_0_2 = 2'h2 == hpOffset ? hpWriteWord_0 : hpFetchLine_0_2; // @[DCache.scala 138:34 DCache.scala 138:34 DCache.scala 137:24]
  wire [31:0] hpWriteLine_0_3 = 2'h3 == hpOffset ? hpWriteWord_0 : hpFetchLine_0_3; // @[DCache.scala 138:34 DCache.scala 138:34 DCache.scala 137:24]
  wire [31:0] _GEN_16 = 2'h1 == hpOffset ? hpFetchLine_1_1 : hpFetchLine_1_0; // @[DCache.scala 135:107 DCache.scala 135:107]
  wire [31:0] _GEN_17 = 2'h2 == hpOffset ? hpFetchLine_1_2 : _GEN_16; // @[DCache.scala 135:107 DCache.scala 135:107]
  wire [31:0] _GEN_18 = 2'h3 == hpOffset ? hpFetchLine_1_3 : _GEN_17; // @[DCache.scala 135:107 DCache.scala 135:107]
  wire [62:0] _GEN_71 = {{31'd0}, _GEN_18}; // @[DCache.scala 135:107]
  wire [62:0] _hpWriteWord_1_T_4 = _hpWriteWord_0_T_3 & _GEN_71; // @[DCache.scala 135:107]
  wire [62:0] _hpWriteWord_1_T_5 = _hpWriteWord_0_T_1 | _hpWriteWord_1_T_4; // @[DCache.scala 135:72]
  wire [31:0] hpWriteWord_1 = _hpWriteWord_1_T_5[31:0]; // @[DCache.scala 130:27 DCache.scala 135:24]
  wire [31:0] hpWriteLine_1_0 = 2'h0 == hpOffset ? hpWriteWord_1 : hpFetchLine_1_0; // @[DCache.scala 138:34 DCache.scala 138:34 DCache.scala 137:24]
  wire [31:0] hpWriteLine_1_1 = 2'h1 == hpOffset ? hpWriteWord_1 : hpFetchLine_1_1; // @[DCache.scala 138:34 DCache.scala 138:34 DCache.scala 137:24]
  wire [31:0] hpWriteLine_1_2 = 2'h2 == hpOffset ? hpWriteWord_1 : hpFetchLine_1_2; // @[DCache.scala 138:34 DCache.scala 138:34 DCache.scala 137:24]
  wire [31:0] hpWriteLine_1_3 = 2'h3 == hpOffset ? hpWriteWord_1 : hpFetchLine_1_3; // @[DCache.scala 138:34 DCache.scala 138:34 DCache.scala 137:24]
  wire [31:0] rdata_0 = meta_1_io_hit ? 32'h0 : hpFetchLine_1_0; // @[DCache.scala 144:21]
  wire [31:0] rdata_1 = meta_1_io_hit ? 32'h0 : hpFetchLine_1_1; // @[DCache.scala 144:21]
  wire [31:0] rdata_2 = meta_1_io_hit ? 32'h0 : hpFetchLine_1_2; // @[DCache.scala 144:21]
  wire [31:0] rdata_3 = meta_1_io_hit ? 32'h0 : hpFetchLine_1_3; // @[DCache.scala 144:21]
  wire [31:0] mpRefillLine_0 = io_bar_resp_bits_rdata[31:0]; // @[DCache.scala 172:56]
  wire [31:0] mpRefillLine_1 = io_bar_resp_bits_rdata[63:32]; // @[DCache.scala 172:56]
  wire [31:0] _GEN_24 = 2'h1 == mpOffset[1:0] ? mpRefillLine_1 : mpRefillLine_0; // @[DCache.scala 146:34 DCache.scala 146:34]
  wire [31:0] mpRefillLine_2 = io_bar_resp_bits_rdata[95:64]; // @[DCache.scala 172:56]
  wire [31:0] _GEN_25 = 2'h2 == mpOffset[1:0] ? mpRefillLine_2 : _GEN_24; // @[DCache.scala 146:34 DCache.scala 146:34]
  wire [31:0] mpRefillLine_3 = io_bar_resp_bits_rdata[127:96]; // @[DCache.scala 172:56]
  wire [31:0] _GEN_26 = 2'h3 == mpOffset[1:0] ? mpRefillLine_3 : _GEN_25; // @[DCache.scala 146:34 DCache.scala 146:34]
  wire [31:0] _GEN_28 = 2'h1 == hpOffset ? rdata_1 : rdata_0; // @[DCache.scala 146:34 DCache.scala 146:34]
  wire [31:0] _GEN_29 = 2'h2 == hpOffset ? rdata_2 : _GEN_28; // @[DCache.scala 146:34 DCache.scala 146:34]
  wire [31:0] _GEN_30 = 2'h3 == hpOffset ? rdata_3 : _GEN_29; // @[DCache.scala 146:34 DCache.scala 146:34]
  wire  _data_0_io_web_T_4 = hpValid & meta_0_io_hit & hpReq_wen; // @[DCache.scala 149:107]
  wire [31:0] _mpWriteWord_T = mpMask & mpReq_wdata; // @[DCache.scala 192:32]
  wire [62:0] _GEN_72 = {{31'd0}, _mpWriteWord_T}; // @[DCache.scala 192:47]
  wire [62:0] _mpWriteWord_T_1 = _GEN_72 << mpShift; // @[DCache.scala 192:47]
  wire [62:0] _GEN_73 = {{31'd0}, mpMask}; // @[DCache.scala 192:81]
  wire [62:0] _mpWriteWord_T_2 = _GEN_73 << mpShift; // @[DCache.scala 192:81]
  wire [62:0] _mpWriteWord_T_3 = ~_mpWriteWord_T_2; // @[DCache.scala 192:72]
  wire [62:0] _GEN_74 = {{31'd0}, _GEN_26}; // @[DCache.scala 192:103]
  wire [62:0] _mpWriteWord_T_5 = _mpWriteWord_T_3 & _GEN_74; // @[DCache.scala 192:103]
  wire [62:0] mpWriteWord = _mpWriteWord_T_1 | _mpWriteWord_T_5; // @[DCache.scala 192:68]
  wire [31:0] mpWriteLine_1 = 2'h1 == mpOffset[1:0] ? mpWriteWord[31:0] : mpRefillLine_1; // @[DCache.scala 194:27 DCache.scala 194:27 DCache.scala 193:17]
  wire [31:0] mpWriteLine_0 = 2'h0 == mpOffset[1:0] ? mpWriteWord[31:0] : mpRefillLine_0; // @[DCache.scala 194:27 DCache.scala 194:27 DCache.scala 193:17]
  wire [31:0] mpWriteLine_3 = 2'h3 == mpOffset[1:0] ? mpWriteWord[31:0] : mpRefillLine_3; // @[DCache.scala 194:27 DCache.scala 194:27 DCache.scala 193:17]
  wire [31:0] mpWriteLine_2 = 2'h2 == mpOffset[1:0] ? mpWriteWord[31:0] : mpRefillLine_2; // @[DCache.scala 194:27 DCache.scala 194:27 DCache.scala 193:17]
  wire [127:0] _data_0_io_dinb_T = {mpWriteLine_3,mpWriteLine_2,mpWriteLine_1,mpWriteLine_0}; // @[DCache.scala 151:74]
  wire [127:0] _data_0_io_dinb_T_1 = mpReq_wen ? _data_0_io_dinb_T : io_bar_resp_bits_rdata; // @[DCache.scala 151:44]
  wire [127:0] _data_0_io_dinb_T_2 = {hpWriteLine_0_3,hpWriteLine_0_2,hpWriteLine_0_1,hpWriteLine_0_0}; // @[DCache.scala 151:133]
  wire  _data_1_io_web_T_4 = hpValid & meta_1_io_hit & hpReq_wen; // @[DCache.scala 149:107]
  wire [127:0] _data_1_io_dinb_T_2 = {hpWriteLine_1_3,hpWriteLine_1_2,hpWriteLine_1_1,hpWriteLine_1_0}; // @[DCache.scala 151:133]
  wire  _meta_0_io_update_T_2 = mpValid ? 1'h0 : _data_0_io_web_T_4; // @[DCache.scala 158:33]
  wire  _meta_1_io_update_T_2 = mpValid ? 1'h0 : _data_1_io_web_T_4; // @[DCache.scala 158:33]
  wire [31:0] _io_bar_req_bits_addr_T_1 = _T_31 ? mpDirtyAddr : mpRefillAddr; // @[DCache.scala 167:46]
  wire [31:0] _mpDirtyAddr_T = {meta_1_io_tagFetch,hpIndex,4'h0}; // @[Cat.scala 30:58]
  wire [127:0] _mpDirtyData_T = {hpFetchLine_1_3,hpFetchLine_1_2,hpFetchLine_1_1,hpFetchLine_1_0}; // @[DCache.scala 185:51]
  wire [31:0] _mpDirtyAddr_T_1 = {meta_0_io_tagFetch,hpIndex,4'h0}; // @[Cat.scala 30:58]
  wire [127:0] _mpDirtyData_T_1 = {hpFetchLine_0_3,hpFetchLine_0_2,hpFetchLine_0_1,hpFetchLine_0_0}; // @[DCache.scala 188:51]
  wire  _GEN_53 = hpTag[0] | _meta_1_io_update_T_2; // @[DCache.scala 202:33 DCache.scala 203:39 DCache.scala 158:27]
  wire  _GEN_54 = hpTag[0] ? _meta_0_io_update_T_2 : 1'h1; // @[DCache.scala 202:33 DCache.scala 158:27 DCache.scala 205:39]
  wire  _GEN_55 = mpState ? _GEN_53 : _meta_1_io_update_T_2; // @[Conditional.scala 39:67 DCache.scala 158:27]
  wire  _GEN_56 = mpState ? _GEN_54 : _meta_0_io_update_T_2; // @[Conditional.scala 39:67 DCache.scala 158:27]
  wire  _GEN_58 = _T_31 | mpState; // @[Conditional.scala 40:58 DCache.scala 199:25 DCache.scala 163:26]
  wire  _GEN_59 = _T_31 ? _meta_1_io_update_T_2 : _GEN_55; // @[Conditional.scala 40:58 DCache.scala 158:27]
  wire  _GEN_60 = _T_31 ? _meta_0_io_update_T_2 : _GEN_56; // @[Conditional.scala 40:58 DCache.scala 158:27]
  DualPortBRAM data_0 ( // @[DCache.scala 54:48]
    .clock(data_0_clock),
    .reset(data_0_reset),
    .io_web(data_0_io_web),
    .io_addra(data_0_io_addra),
    .io_addrb(data_0_io_addrb),
    .io_dinb(data_0_io_dinb),
    .io_douta(data_0_io_douta)
  );
  DualPortBRAM data_1 ( // @[DCache.scala 54:48]
    .clock(data_1_clock),
    .reset(data_1_reset),
    .io_web(data_1_io_web),
    .io_addra(data_1_io_addra),
    .io_addrb(data_1_io_addrb),
    .io_dinb(data_1_io_dinb),
    .io_douta(data_1_io_douta)
  );
  MetaDataBRAM meta_0 ( // @[DCache.scala 55:48]
    .clock(meta_0_clock),
    .reset(meta_0_reset),
    .io_indexFetch(meta_0_io_indexFetch),
    .io_indexUpdate(meta_0_io_indexUpdate),
    .io_tagUpdate(meta_0_io_tagUpdate),
    .io_update(meta_0_io_update),
    .io_write(meta_0_io_write),
    .io_hit(meta_0_io_hit),
    .io_tagFetch(meta_0_io_tagFetch)
  );
  MetaDataBRAM meta_1 ( // @[DCache.scala 55:48]
    .clock(meta_1_clock),
    .reset(meta_1_reset),
    .io_indexFetch(meta_1_io_indexFetch),
    .io_indexUpdate(meta_1_io_indexUpdate),
    .io_tagUpdate(meta_1_io_tagUpdate),
    .io_update(meta_1_io_update),
    .io_write(meta_1_io_write),
    .io_hit(meta_1_io_hit),
    .io_tagFetch(meta_1_io_tagFetch)
  );
  assign io_cpu_req_ready = io_cpu_resp_valid; // @[DCache.scala 173:22]
  assign io_cpu_resp_valid = hpRespValid | mpRespValid; // @[DCache.scala 141:43]
  assign io_cpu_resp_bits_rdata = mpValid ? _GEN_26 : _GEN_30; // @[DCache.scala 146:34]
  assign io_bar_req_bits_addr = mpValid ? _io_bar_req_bits_addr_T_1 : io_cpu_req_bits_addr; // @[DCache.scala 167:33]
  assign io_bar_req_bits_wen = mpValid ? _T_31 : io_cpu_req_bits_wen; // @[DCache.scala 170:33]
  assign io_bar_req_bits_wdata = mpValid ? mpDirtyData : {{96'd0}, io_cpu_req_bits_wdata}; // @[DCache.scala 168:33]
  assign io_bar_req_bits_mtype = io_cpu_req_bits_mtype; // @[DCache.scala 169:27]
  assign io_dbg_hit = meta_0_io_hit | meta_1_io_hit; // @[DCache.scala 109:31]
  assign io_dbg_hitWay = _hpRespValid_T & meta_1_io_hit; // @[DCache.scala 114:33]
  assign io_dbg_replaceWay = hpTag[0]; // @[DCache.scala 115:31]
  assign data_0_clock = clock;
  assign data_0_reset = reset;
  assign data_0_io_web = mpValid ? ~mpTag[0] & mpWriteCache : hpValid & meta_0_io_hit & hpReq_wen; // @[DCache.scala 149:30]
  assign data_0_io_addra = io_cpu_req_bits_addr[11:4]; // @[DCache.scala 65:40]
  assign data_0_io_addrb = mpValid ? mpIndex : hpIndex; // @[DCache.scala 150:32]
  assign data_0_io_dinb = mpValid ? _data_0_io_dinb_T_1 : _data_0_io_dinb_T_2; // @[DCache.scala 151:31]
  assign data_1_clock = clock;
  assign data_1_reset = reset;
  assign data_1_io_web = mpValid ? mpTag[0] & mpWriteCache : hpValid & meta_1_io_hit & hpReq_wen; // @[DCache.scala 149:30]
  assign data_1_io_addra = io_cpu_req_bits_addr[11:4]; // @[DCache.scala 65:40]
  assign data_1_io_addrb = mpValid ? mpIndex : hpIndex; // @[DCache.scala 150:32]
  assign data_1_io_dinb = mpValid ? _data_0_io_dinb_T_1 : _data_1_io_dinb_T_2; // @[DCache.scala 151:31]
  assign meta_0_clock = clock;
  assign meta_0_reset = reset;
  assign meta_0_io_indexFetch = io_cpu_req_bits_addr[11:4]; // @[DCache.scala 65:40]
  assign meta_0_io_indexUpdate = mpValid ? mpIndex : hpIndex; // @[DCache.scala 155:38]
  assign meta_0_io_tagUpdate = mpValid ? mpTag : hpTag; // @[DCache.scala 156:38]
  assign meta_0_io_update = mpValid ? _GEN_60 : _meta_0_io_update_T_2; // @[DCache.scala 196:20 DCache.scala 158:27]
  assign meta_0_io_write = mpValid ? mpReq_wen : hpReq_wen; // @[DCache.scala 157:33]
  assign meta_1_clock = clock;
  assign meta_1_reset = reset;
  assign meta_1_io_indexFetch = io_cpu_req_bits_addr[11:4]; // @[DCache.scala 65:40]
  assign meta_1_io_indexUpdate = mpValid ? mpIndex : hpIndex; // @[DCache.scala 155:38]
  assign meta_1_io_tagUpdate = mpValid ? mpTag : hpTag; // @[DCache.scala 156:38]
  assign meta_1_io_update = mpValid ? _GEN_59 : _meta_1_io_update_T_2; // @[DCache.scala 196:20 DCache.scala 158:27]
  assign meta_1_io_write = mpValid ? mpReq_wen : hpReq_wen; // @[DCache.scala 157:33]
  always @(posedge clock) begin
    if (reset) begin // @[DCache.scala 85:26]
      mpValid <= 1'h0; // @[DCache.scala 85:26]
    end else if (_hpReq_T) begin // @[DCache.scala 175:21]
      mpValid <= _hpValid_T_1; // @[DCache.scala 176:21]
    end
    if (reset) begin // @[DCache.scala 163:26]
      mpState <= 1'h0; // @[DCache.scala 163:26]
    end else if (mpValid) begin // @[DCache.scala 196:20]
      mpState <= _GEN_58;
    end
    if (_hpReq_T) begin // @[Reg.scala 16:19]
      hpReq_addr <= io_cpu_req_bits_addr; // @[Reg.scala 16:23]
    end
    if (_hpReq_T) begin // @[Reg.scala 16:19]
      hpReq_wen <= io_cpu_req_bits_wen; // @[Reg.scala 16:23]
    end
    if (_hpReq_T) begin // @[Reg.scala 16:19]
      hpReq_wdata <= io_cpu_req_bits_wdata; // @[Reg.scala 16:23]
    end
    if (_hpReq_T) begin // @[Reg.scala 16:19]
      hpReq_mtype <= io_cpu_req_bits_mtype; // @[Reg.scala 16:23]
    end
    if (_hpReq_T) begin // @[Reg.scala 16:19]
      hpIndex <= arIndex; // @[Reg.scala 16:23]
    end
    if (_hpReq_T) begin // @[Reg.scala 16:19]
      hpTag <= arTag; // @[Reg.scala 16:23]
    end
    if (_hpReq_T) begin // @[Reg.scala 16:19]
      hpOffset <= arOffset; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[DCache.scala 79:30]
      hpValid <= 1'h0; // @[DCache.scala 79:30]
    end else if (hpValid & ~_hpRespValid_T | mpStall) begin // @[DCache.scala 111:19]
      hpValid <= 1'h0;
    end else begin
      hpValid <= io_cpu_req_valid;
    end
    if (reset) begin // @[DCache.scala 83:26]
      mpReq_wen <= 1'h0; // @[DCache.scala 83:26]
    end else if (_hpReq_T) begin // @[DCache.scala 175:21]
      mpReq_wen <= hpReq_wen; // @[DCache.scala 177:21]
    end
    if (reset) begin // @[DCache.scala 83:26]
      mpReq_wdata <= 32'h0; // @[DCache.scala 83:26]
    end else if (_hpReq_T) begin // @[DCache.scala 175:21]
      mpReq_wdata <= hpReq_wdata; // @[DCache.scala 177:21]
    end
    if (_hpReq_T) begin // @[DCache.scala 175:21]
      if (hpTag[0]) begin // @[DCache.scala 183:25]
        mpDirtyAddr <= _mpDirtyAddr_T; // @[DCache.scala 184:25]
      end else begin
        mpDirtyAddr <= _mpDirtyAddr_T_1; // @[DCache.scala 187:25]
      end
    end
    if (_hpReq_T) begin // @[DCache.scala 175:21]
      if (hpTag[0]) begin // @[DCache.scala 183:25]
        mpDirtyData <= _mpDirtyData_T; // @[DCache.scala 185:25]
      end else begin
        mpDirtyData <= _mpDirtyData_T_1; // @[DCache.scala 188:25]
      end
    end
    if (reset) begin // @[DCache.scala 93:27]
      mpOffset <= 4'h0; // @[DCache.scala 93:27]
    end else if (_hpReq_T) begin // @[DCache.scala 175:21]
      mpOffset <= {{2'd0}, hpOffset}; // @[DCache.scala 180:21]
    end
    if (reset) begin // @[DCache.scala 94:27]
      mpIndex <= 8'h0; // @[DCache.scala 94:27]
    end else if (_hpReq_T) begin // @[DCache.scala 175:21]
      mpIndex <= hpIndex; // @[DCache.scala 178:21]
    end
    if (reset) begin // @[DCache.scala 95:27]
      mpTag <= 20'h0; // @[DCache.scala 95:27]
    end else if (_hpReq_T) begin // @[DCache.scala 175:21]
      mpTag <= hpTag; // @[DCache.scala 179:21]
    end
    if (_hpReq_T) begin // @[DCache.scala 175:21]
      if (2'h1 == hpReq_mtype) begin // @[Mux.scala 80:57]
        mpMask <= 32'hffff;
      end else if (2'h0 == hpReq_mtype) begin // @[Mux.scala 80:57]
        mpMask <= 32'hff;
      end else begin
        mpMask <= 32'hffffffff;
      end
    end
    if (_hpReq_T) begin // @[DCache.scala 175:21]
      mpShift <= hpShift; // @[DCache.scala 182:21]
    end
    REG <= data_0_io_web & data_0_io_addra == data_0_io_addrb; // @[DCache.scala 118:54]
    REG_1_0 <= _WIRE_1[31:0]; // @[DCache.scala 119:65]
    REG_1_1 <= _WIRE_1[63:32]; // @[DCache.scala 119:65]
    REG_1_2 <= _WIRE_1[95:64]; // @[DCache.scala 119:65]
    REG_1_3 <= _WIRE_1[127:96]; // @[DCache.scala 119:65]
    REG_2 <= data_1_io_web & data_1_io_addra == data_1_io_addrb; // @[DCache.scala 118:54]
    REG_3_0 <= _WIRE_5[31:0]; // @[DCache.scala 119:65]
    REG_3_1 <= _WIRE_5[63:32]; // @[DCache.scala 119:65]
    REG_3_2 <= _WIRE_5[95:64]; // @[DCache.scala 119:65]
    REG_3_3 <= _WIRE_5[127:96]; // @[DCache.scala 119:65]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mpValid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  mpState = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  hpReq_addr = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  hpReq_wen = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  hpReq_wdata = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  hpReq_mtype = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  hpIndex = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  hpTag = _RAND_7[19:0];
  _RAND_8 = {1{`RANDOM}};
  hpOffset = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  hpValid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  mpReq_wen = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  mpReq_wdata = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  mpDirtyAddr = _RAND_12[31:0];
  _RAND_13 = {4{`RANDOM}};
  mpDirtyData = _RAND_13[127:0];
  _RAND_14 = {1{`RANDOM}};
  mpOffset = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  mpIndex = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  mpTag = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  mpMask = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  mpShift = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  REG = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  REG_1_0 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  REG_1_1 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  REG_1_2 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  REG_1_3 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  REG_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  REG_3_0 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  REG_3_1 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  REG_3_2 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  REG_3_3 = _RAND_28[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Test(
  input         clock,
  input         reset,
  output        io_dbg_hit,
  output        io_dbg_hitWay,
  output        io_dbg_replaceWay,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input         io_cpu_req_bits_wen,
  input  [31:0] io_cpu_req_bits_wdata,
  input  [1:0]  io_cpu_req_bits_mtype,
  input         io_cpu_resp_ready,
  output        io_cpu_resp_valid,
  output [31:0] io_cpu_resp_bits_rdata
);
  wire  dcache_clock; // @[Test.scala 36:24]
  wire  dcache_reset; // @[Test.scala 36:24]
  wire  dcache_io_cpu_req_ready; // @[Test.scala 36:24]
  wire  dcache_io_cpu_req_valid; // @[Test.scala 36:24]
  wire [31:0] dcache_io_cpu_req_bits_addr; // @[Test.scala 36:24]
  wire  dcache_io_cpu_req_bits_wen; // @[Test.scala 36:24]
  wire [31:0] dcache_io_cpu_req_bits_wdata; // @[Test.scala 36:24]
  wire [1:0] dcache_io_cpu_req_bits_mtype; // @[Test.scala 36:24]
  wire  dcache_io_cpu_resp_valid; // @[Test.scala 36:24]
  wire [31:0] dcache_io_cpu_resp_bits_rdata; // @[Test.scala 36:24]
  wire [31:0] dcache_io_bar_req_bits_addr; // @[Test.scala 36:24]
  wire  dcache_io_bar_req_bits_wen; // @[Test.scala 36:24]
  wire [127:0] dcache_io_bar_req_bits_wdata; // @[Test.scala 36:24]
  wire [1:0] dcache_io_bar_req_bits_mtype; // @[Test.scala 36:24]
  wire [127:0] dcache_io_bar_resp_bits_rdata; // @[Test.scala 36:24]
  wire  dcache_io_dbg_hit; // @[Test.scala 36:24]
  wire  dcache_io_dbg_hitWay; // @[Test.scala 36:24]
  wire  dcache_io_dbg_replaceWay; // @[Test.scala 36:24]
  wire  dmem_clka; // @[Test.scala 37:24]
  wire [31:0] dmem_addra; // @[Test.scala 37:24]
  wire [31:0] dmem_dina; // @[Test.scala 37:24]
  wire  dmem_wea; // @[Test.scala 37:24]
  wire [31:0] dmem_douta; // @[Test.scala 37:24]
  wire [1:0] dmem_mtype; // @[Test.scala 37:24]
  DCache dcache ( // @[Test.scala 36:24]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_cpu_req_ready(dcache_io_cpu_req_ready),
    .io_cpu_req_valid(dcache_io_cpu_req_valid),
    .io_cpu_req_bits_addr(dcache_io_cpu_req_bits_addr),
    .io_cpu_req_bits_wen(dcache_io_cpu_req_bits_wen),
    .io_cpu_req_bits_wdata(dcache_io_cpu_req_bits_wdata),
    .io_cpu_req_bits_mtype(dcache_io_cpu_req_bits_mtype),
    .io_cpu_resp_valid(dcache_io_cpu_resp_valid),
    .io_cpu_resp_bits_rdata(dcache_io_cpu_resp_bits_rdata),
    .io_bar_req_bits_addr(dcache_io_bar_req_bits_addr),
    .io_bar_req_bits_wen(dcache_io_bar_req_bits_wen),
    .io_bar_req_bits_wdata(dcache_io_bar_req_bits_wdata),
    .io_bar_req_bits_mtype(dcache_io_bar_req_bits_mtype),
    .io_bar_resp_bits_rdata(dcache_io_bar_resp_bits_rdata),
    .io_dbg_hit(dcache_io_dbg_hit),
    .io_dbg_hitWay(dcache_io_dbg_hitWay),
    .io_dbg_replaceWay(dcache_io_dbg_replaceWay)
  );
  RAM_B dmem ( // @[Test.scala 37:24]
    .clka(dmem_clka),
    .addra(dmem_addra),
    .dina(dmem_dina),
    .wea(dmem_wea),
    .douta(dmem_douta),
    .mtype(dmem_mtype)
  );
  assign io_dbg_hit = dcache_io_dbg_hit; // @[Test.scala 49:19]
  assign io_dbg_hitWay = dcache_io_dbg_hitWay; // @[Test.scala 49:19]
  assign io_dbg_replaceWay = dcache_io_dbg_replaceWay; // @[Test.scala 49:19]
  assign io_cpu_req_ready = dcache_io_cpu_req_ready; // @[Test.scala 48:19]
  assign io_cpu_resp_valid = dcache_io_cpu_resp_valid; // @[Test.scala 48:19]
  assign io_cpu_resp_bits_rdata = dcache_io_cpu_resp_bits_rdata; // @[Test.scala 48:19]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_cpu_req_valid = io_cpu_req_valid; // @[Test.scala 48:19]
  assign dcache_io_cpu_req_bits_addr = io_cpu_req_bits_addr; // @[Test.scala 48:19]
  assign dcache_io_cpu_req_bits_wen = io_cpu_req_bits_wen; // @[Test.scala 48:19]
  assign dcache_io_cpu_req_bits_wdata = io_cpu_req_bits_wdata; // @[Test.scala 48:19]
  assign dcache_io_cpu_req_bits_mtype = io_cpu_req_bits_mtype; // @[Test.scala 48:19]
  assign dcache_io_bar_resp_bits_rdata = {{96'd0}, dmem_douta}; // @[Test.scala 43:35]
  assign dmem_clka = clock; // @[Test.scala 38:19]
  assign dmem_addra = dcache_io_bar_req_bits_addr; // @[Test.scala 41:19]
  assign dmem_dina = dcache_io_bar_req_bits_wdata[31:0]; // @[Test.scala 42:19]
  assign dmem_wea = dcache_io_bar_req_bits_wen; // @[Test.scala 40:19]
  assign dmem_mtype = dcache_io_bar_req_bits_mtype; // @[Test.scala 39:19]
endmodule
//-------------------------------------
module RAM_B(
    input [31:0] addra,
    input clka,      // normal clock
    input[127:0] dina,
    input wea, 
    output[127:0] douta,
    input[1:0] mtype
);

    reg[7:0] data[0:511];

    initial	begin
        $readmemh("ram.hex", data);
    end

    always @(posedge clka) begin
        if (wea & ~|addra[30:9]) begin
            data[addra[8:0] + 15] <= dina[127 : 120];
            data[addra[8:0] + 14] <= dina[119 : 112];
            data[addra[8:0] + 13] <= dina[111 : 104];
            data[addra[8:0] + 12] <= dina[103 : 96];
            data[addra[8:0] + 11] <= dina[95  : 88];
            data[addra[8:0] + 10] <= dina[87  : 80];
            data[addra[8:0] + 9]  <= dina[79  : 72];
            data[addra[8:0] + 8]  <= dina[71  : 64];
            data[addra[8:0] + 7]  <= dina[63  : 56];
            data[addra[8:0] + 6]  <= dina[55  : 48];
            data[addra[8:0] + 5]  <= dina[47  : 40];
            data[addra[8:0] + 4]  <= dina[39  : 32];
            data[addra[8:0] + 3]  <= dina[31  : 24];
            data[addra[8:0] + 2]  <= dina[23  : 16];
            data[addra[8:0] + 1]  <= dina[15  : 8];
            data[addra[8:0]]      <= dina[7   : 0];
        end
    end
    
    assign douta = addra[30:9] ? 128'b0 :
                   {data[addra[8:0] + 15],
                    data[addra[8:0] + 14],
                    data[addra[8:0] + 13],
                    data[addra[8:0] + 12],
                    data[addra[8:0] + 11], 
                    data[addra[8:0] + 10], 
                    data[addra[8:0] + 9], 
                    data[addra[8:0] + 8],
                    data[addra[8:0] + 7],
                    data[addra[8:0] + 6],
                    data[addra[8:0] + 5],
                    data[addra[8:0] + 4],
                    data[addra[8:0] + 3], 
                    data[addra[8:0] + 2], 
                    data[addra[8:0] + 1], 
                    data[addra[8:0]]};

endmodule